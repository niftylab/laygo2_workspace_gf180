* NGSPICE file created from dec3to8.ext - technology: gf180mcuC

.subckt dec3to8 A0 A1 A2 EN Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 VDD VSS
X0 and4_5.nand0.OUT A0 a_20460_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1 and4_5.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2 a_15420_1092# and4_3.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3 and4_4.nand1.OUT and4_5.nand1.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4 Y1 and4_1.nand1.OUT a_8220_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5 VDD A0 and4_5.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6 and4_0.nand0.OUT and4_6.nand0.A a_2460_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7 Y3 and4_3.nand1.OUT a_15420_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8 a_17940_306# A2 and4_4.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9 and4_1.nand1.OUT and4_5.nand1.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10 VSS and4_3.nand0.OUT Y3 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11 Y2 and4_2.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12 and4_7.nand1.OUT A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X13 VSS A0 and4_6.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X14 and4_3.nand1.OUT and4_3.nand1.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X15 Y6 and4_6.nand1.OUT a_26220_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X16 a_16860_306# and4_6.nand0.A and4_4.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X17 a_25140_306# A2 and4_6.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X18 VSS A1 a_14340_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X19 VSS and4_5.nand0.OUT Y5 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X20 VSS EN a_13260_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X21 and4_0.nand1.OUT and4_3.nand1.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X22 VDD and4_3.nand0.OUT a_15420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X23 and4_6.nand1.OUT A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X24 a_24060_306# and4_6.nand0.A and4_6.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X25 and4_1.nand0.OUT A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X26 VSS and4_5.nand1.B a_21540_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X27 and4_2.nand1.OUT A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X28 and4_4.nand1.OUT A2 a_17940_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X29 and4_6.nand0.A A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X30 Y3 and4_3.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X31 a_7140_306# and4_3.nand1.A and4_1.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X32 a_15420_1092# and4_3.nand1.OUT Y3 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X33 and4_6.nand0.A A0 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X34 VSS EN a_20460_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X35 VSS and4_0.nand0.OUT Y0 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X36 VDD and4_5.nand1.B and4_1.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X37 and4_4.nand0.OUT and4_6.nand0.A a_16860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X38 VDD EN and4_2.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X39 VDD A2 and4_7.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X40 and4_6.nand1.OUT A2 a_25140_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X41 a_14340_306# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X42 and4_5.nand1.OUT A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X43 Y5 and4_5.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X44 a_6060_306# A0 and4_1.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X45 and4_6.nand0.OUT and4_6.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X46 VSS and4_5.nand1.B a_3540_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X47 VSS A2 and4_3.nand1.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X48 VSS and4_3.nand1.OUT Y3 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X49 a_27660_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X50 and4_6.nand0.OUT and4_6.nand0.A a_24060_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X51 a_21540_306# and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X52 VSS EN a_2460_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X53 and4_3.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X54 VDD A1 and4_6.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X55 VDD and4_3.nand1.A and4_0.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X56 VDD A0 and4_1.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X57 VDD EN and4_7.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X58 VSS and4_5.nand1.OUT Y5 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X59 and4_1.nand1.OUT and4_3.nand1.A a_7140_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X60 VDD A1 and4_2.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X61 Y0 and4_0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X62 VDD A0 and4_6.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X63 a_9660_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X64 and4_1.nand0.OUT A0 a_6060_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X65 a_19020_1092# and4_4.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X66 VSS and4_7.nand1.OUT Y7 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X67 VSS and4_4.nand0.OUT Y4 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X68 a_3540_306# and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X69 Y3 and4_3.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X70 VDD EN and4_0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X71 and4_3.nand1.A A2 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X72 VDD A2 and4_5.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X73 VDD and4_6.nand0.A and4_6.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X74 VSS and4_0.nand1.OUT Y0 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X75 VSS and4_5.nand1.B a_17940_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X76 Y4 and4_4.nand1.OUT a_19020_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X77 a_28740_306# A2 and4_7.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X78 a_8220_1092# and4_1.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X79 VSS and4_6.nand0.OUT Y6 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X80 Y5 and4_5.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X81 a_27660_306# A0 and4_7.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X82 VSS A1 a_25140_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X83 a_10740_306# and4_3.nand1.A and4_2.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X84 VDD EN and4_5.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X85 Y7 and4_7.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X86 a_26220_1092# and4_6.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X87 VSS EN a_24060_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X88 a_9660_306# and4_6.nand0.A and4_2.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X89 VSS and4_1.nand0.OUT Y1 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X90 and4_7.nand1.OUT A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X91 Y0 and4_0.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X92 and4_1.nand1.OUT and4_3.nand1.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X93 a_11820_1092# and4_2.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X94 and4_7.nand1.OUT A2 a_28740_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X95 Y6 and4_6.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X96 VSS and4_5.nand1.B a_7140_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X97 and4_4.nand0.OUT and4_6.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X98 VDD and4_1.nand0.OUT a_8220_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X99 a_19020_1092# and4_4.nand1.OUT Y4 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X100 and4_7.nand0.OUT A0 a_27660_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X101 and4_2.nand1.OUT and4_3.nand1.A a_10740_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X102 Y2 and4_2.nand1.OUT a_11820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X103 a_25140_306# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X104 VSS EN a_6060_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X105 and4_0.nand1.OUT and4_5.nand1.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X106 and4_6.nand1.OUT A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X107 VDD and4_5.nand1.B and4_4.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X108 VSS and4_6.nand1.OUT Y6 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X109 a_13260_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X110 and4_2.nand0.OUT and4_6.nand0.A a_9660_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X111 and4_5.nand1.B A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X112 a_8220_1092# and4_1.nand1.OUT Y1 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X113 Y1 and4_1.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X114 and4_4.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X115 VDD and4_6.nand0.OUT a_26220_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X116 VDD A1 and4_7.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X117 a_7140_306# and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X118 VDD and4_3.nand1.A and4_1.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X119 a_20460_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X120 VDD and4_2.nand0.OUT a_11820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X121 and4_5.nand1.OUT and4_5.nand1.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X122 and4_0.nand0.OUT and4_6.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X123 VSS and4_1.nand1.OUT Y1 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X124 VDD and4_3.nand1.A and4_3.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X125 VDD and4_6.nand0.A and4_4.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X126 a_26220_1092# and4_6.nand1.OUT Y6 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X127 and4_1.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X128 and4_2.nand0.OUT and4_6.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X129 a_11820_1092# and4_2.nand1.OUT Y2 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X130 VDD A1 and4_5.nand1.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X131 VDD and4_5.nand1.B and4_0.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X132 VDD A2 and4_6.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X133 a_2460_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X134 Y7 and4_7.nand1.OUT a_29820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X135 a_14340_306# and4_3.nand1.A and4_3.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X136 and4_5.nand0.OUT A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X137 VDD EN and4_3.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X138 VSS EN a_16860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X139 and4_6.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X140 a_21540_306# A2 and4_5.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X141 VDD and4_5.nand1.B and4_5.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X142 Y4 and4_4.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X143 a_20460_306# A0 and4_5.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X144 a_29820_1092# and4_7.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X145 a_17940_306# and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X146 VDD and4_6.nand0.A and4_2.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X147 VSS and4_4.nand1.OUT Y4 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X148 a_3540_306# and4_3.nand1.A and4_0.nand1.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X149 and4_5.nand1.B A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X150 VSS A1 and4_5.nand1.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X151 and4_4.nand1.OUT A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X152 a_29820_1092# and4_7.nand1.OUT Y7 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X153 and4_5.nand1.OUT A2 a_21540_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X154 a_2460_306# and4_6.nand0.A and4_0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X155 a_4620_1092# and4_0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X156 VDD and4_4.nand0.OUT a_19020_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X157 a_24060_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X158 and4_3.nand1.OUT A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X159 Y0 and4_0.nand1.OUT a_4620_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X160 VDD and4_7.nand0.OUT a_29820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X161 Y4 and4_4.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X162 and4_0.nand1.OUT and4_3.nand1.A a_3540_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X163 and4_3.nand1.A A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X164 a_22620_1092# and4_5.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X165 VSS and4_7.nand0.OUT Y7 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X166 a_6060_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X167 VDD A2 and4_4.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X168 and4_7.nand0.OUT A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X169 Y6 and4_6.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X170 and4_2.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X171 and4_2.nand1.OUT and4_3.nand1.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X172 and4_3.nand0.OUT A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X173 Y5 and4_5.nand1.OUT a_22620_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X174 VDD and4_0.nand0.OUT a_4620_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X175 VSS A1 a_28740_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X176 VSS and4_2.nand0.OUT Y2 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X177 VDD A1 and4_3.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X178 VSS EN a_27660_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X179 a_13260_306# A0 and4_3.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X180 a_4620_1092# and4_0.nand1.OUT Y0 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X181 VDD EN and4_4.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X182 VSS A1 a_10740_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X183 Y1 and4_1.nand1.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X184 and4_7.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X185 VDD A2 and4_3.nand1.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X186 VDD and4_5.nand0.OUT a_22620_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X187 Y7 and4_7.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X188 VDD EN and4_1.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X189 VDD A0 and4_7.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X190 a_28740_306# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X191 and4_3.nand1.OUT and4_3.nand1.A a_14340_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X192 Y2 and4_2.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X193 VSS EN a_9660_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X194 VDD and4_3.nand1.A and4_2.nand1.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X195 a_22620_1092# and4_5.nand1.OUT Y5 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X196 and4_0.nand0.OUT EN VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X197 VDD A0 and4_3.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X198 a_16860_306# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X199 and4_3.nand0.OUT A0 a_13260_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X200 a_10740_306# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X201 VDD EN and4_6.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X202 VDD and4_6.nand0.A and4_0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X203 VSS and4_2.nand1.OUT Y2 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
.ends

