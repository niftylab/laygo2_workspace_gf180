magic
tech gf180mcuC
magscale 1 10
timestamp 1684124021
<< metal2 >>
rect -105 -28 -91 28
rect 91 -28 105 28
<< via2 >>
rect -91 -28 91 28
<< metal3 >>
rect -105 -28 -91 28
rect 91 -28 105 28
<< end >>
