magic
tech gf180mcuC
magscale 1 10
timestamp 1683428588
<< nmos >>
rect 60 306 120 476
rect 240 306 300 476
<< ndiff >>
rect -60 459 60 476
rect -60 413 -30 459
rect 30 413 60 459
rect -60 365 60 413
rect -60 319 -30 365
rect 30 319 60 365
rect -60 306 60 319
rect 120 459 240 476
rect 120 413 150 459
rect 210 413 240 459
rect 120 365 240 413
rect 120 319 150 365
rect 210 319 240 365
rect 120 306 240 319
rect 300 459 420 476
rect 300 413 330 459
rect 390 413 420 459
rect 300 365 420 413
rect 300 319 330 365
rect 390 319 420 365
rect 300 306 420 319
<< ndiffc >>
rect -30 413 30 459
rect -30 319 30 365
rect 150 413 210 459
rect 150 319 210 365
rect 330 413 390 459
rect 330 319 390 365
<< polysilicon >>
rect -44 650 120 666
rect -44 580 -30 650
rect 30 580 120 650
rect -44 566 120 580
rect 60 476 120 566
rect 240 650 404 666
rect 240 580 330 650
rect 390 580 404 650
rect 240 566 404 580
rect 240 476 300 566
rect 60 262 120 306
rect 240 262 300 306
<< polycontact >>
rect -30 580 30 650
rect 330 580 390 650
<< metal1 >>
rect -44 650 44 672
rect -44 580 -30 650
rect 30 580 44 650
rect -44 560 44 580
rect 316 650 404 672
rect 316 580 330 650
rect 390 580 404 650
rect 316 560 404 580
rect -44 459 44 476
rect -44 413 -30 459
rect 30 413 44 459
rect -44 365 44 413
rect -44 319 -30 365
rect 30 319 44 365
rect -44 280 44 319
rect 136 459 224 476
rect 136 413 150 459
rect 210 413 224 459
rect 136 365 224 413
rect 136 319 150 365
rect 210 319 224 365
rect 136 280 224 319
rect 316 459 404 476
rect 316 413 330 459
rect 390 413 404 459
rect 316 365 404 413
rect 316 319 330 365
rect 390 319 404 365
rect 316 280 404 319
<< end >>
