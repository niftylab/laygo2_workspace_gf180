magic
tech gf180mcuC
timestamp 1683993426
<< properties >>
string FIXED_BBOX 0 0 18 78
<< end >>
