magic
tech gf180mcuC
magscale 1 5
timestamp 1683702384
<< metal1 >>
rect -22 13 22 14
rect -22 -13 -15 13
rect 15 -13 22 13
rect -22 -14 22 -13
<< via1 >>
rect -15 -13 15 13
<< metal2 >>
rect -22 13 22 14
rect -22 -13 -15 13
rect 15 -13 22 13
rect -22 -14 22 -13
<< end >>
