magic
tech gf180mcuC
magscale 1 10
timestamp 1684136783
<< nwell >>
rect -180 -90 540 570
<< pmos >>
rect 60 136 120 476
rect 240 136 300 476
<< pdiff >>
rect -60 450 60 476
rect -60 390 -31 450
rect 31 390 60 450
rect -60 330 60 390
rect -60 270 -31 330
rect 31 270 60 330
rect -60 210 60 270
rect -60 150 -31 210
rect 31 150 60 210
rect -60 136 60 150
rect 120 450 240 476
rect 120 390 149 450
rect 211 390 240 450
rect 120 330 240 390
rect 120 270 149 330
rect 211 270 240 330
rect 120 210 240 270
rect 120 150 149 210
rect 211 150 240 210
rect 120 136 240 150
rect 300 450 420 476
rect 300 390 329 450
rect 391 390 420 450
rect 300 330 420 390
rect 300 270 329 330
rect 391 270 420 330
rect 300 210 420 270
rect 300 150 329 210
rect 391 150 420 210
rect 300 136 420 150
<< pdiffc >>
rect -31 390 31 450
rect -31 270 31 330
rect -31 150 31 210
rect 149 390 211 450
rect 149 270 211 330
rect 149 150 211 210
rect 329 390 391 450
rect 329 270 391 330
rect 329 150 391 210
<< nsubdiff >>
rect -40 55 40 70
rect -40 -45 -25 55
rect 25 -45 40 55
rect -40 -60 40 -45
rect 320 55 400 70
rect 320 -45 335 55
rect 385 -45 400 55
rect 320 -60 400 -45
<< nsubdiffcont >>
rect -25 -45 25 55
rect 335 -45 385 55
<< polysilicon >>
rect 60 650 300 666
rect 60 580 150 650
rect 210 580 300 650
rect 60 566 300 580
rect 60 476 120 566
rect 240 476 300 566
rect 60 84 120 136
rect 240 84 300 136
<< polycontact >>
rect 150 580 210 650
<< metal1 >>
rect 136 650 224 672
rect 136 580 150 650
rect 210 580 224 650
rect 136 560 224 580
rect -44 450 44 476
rect -44 390 -31 450
rect 31 390 44 450
rect -44 330 44 390
rect -44 270 -31 330
rect 31 270 44 330
rect -44 210 44 270
rect -44 150 -31 210
rect 31 150 44 210
rect -44 136 44 150
rect 136 450 224 476
rect 136 390 149 450
rect 211 390 224 450
rect 136 330 224 390
rect 136 270 149 330
rect 211 270 224 330
rect 136 210 224 270
rect 136 150 149 210
rect 211 150 224 210
rect 136 136 224 150
rect 316 450 404 476
rect 316 390 329 450
rect 391 390 404 450
rect 316 330 404 390
rect 316 270 329 330
rect 391 270 404 330
rect 316 210 404 270
rect 316 150 329 210
rect 391 150 404 210
rect 316 136 404 150
rect -44 74 44 84
rect -44 -74 -30 74
rect 30 -74 44 74
rect -44 -84 44 -74
rect 316 74 404 84
rect 316 -74 330 74
rect 390 -74 404 74
rect 316 -84 404 -74
<< via1 >>
rect -30 55 30 74
rect -30 -45 -25 55
rect -25 -45 25 55
rect 25 -45 30 55
rect -30 -74 30 -45
rect 330 55 390 74
rect 330 -45 335 55
rect 335 -45 385 55
rect 385 -45 390 55
rect 330 -74 390 -45
<< metal2 >>
rect -50 74 50 84
rect -50 -74 -30 74
rect 30 -74 50 74
rect -50 -84 50 -74
rect 310 74 410 84
rect 310 -74 330 74
rect 390 -74 410 74
rect 310 -84 410 -74
<< end >>
