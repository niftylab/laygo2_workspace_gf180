* NGSPICE file created from dff_byte_right.ext - technology: gf180mcuC

.subckt dff_byte_right CLK Di<0> Di<1> Di<2> Di<3> Di<4> Di<5> Di<6> Di<7> Do<0> Do<1>
+ Do<2> Do<3> Do<4> Do<5> Do<6> Do<7> RE SEL WE VSS VDD
X0 VSS a_17860_140# a_17760_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1 Do<2> tinv7.EN a_20460_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2 a_22620_680# a_22410_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3 VSS a_35760_190# a_36420_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4 VDD a_15420_680# a_15380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5 dff_2.O tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6 a_15380_190# a_14590_140# a_15210_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7 a_20460_1092# tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8 VDD tinv6.I a_34860_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9 a_18190_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10 a_14820_190# dff_7.CLK a_14260_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11 VSS a_19020_680# tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12 dff_6.O tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X13 VDD a_21360_190# a_22020_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X14 VDD RE tinv7.ENB VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X15 dff_5.O tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X16 a_29820_680# a_29610_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X17 a_22580_190# a_21790_140# a_22410_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X18 a_14260_140# dff_7.CLK a_14490_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X19 a_20460_1092# tinv7.ENB Do<2> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X20 VDD a_25060_140# a_24960_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X21 cgate0.latch0.I2.I cgate0.latch0.I1.ENB a_2460_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X22 a_22020_190# dff_7.CLK a_21460_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X23 VDD a_32160_190# a_32820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X24 a_11500_1090# a_10560_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X25 VDD cgate0.nand0.OUT dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X26 VDD a_10660_140# a_10560_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X27 a_18420_1090# a_18190_140# a_17860_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X28 a_15420_680# a_15210_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X29 a_17860_140# a_18190_140# a_18090_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X30 a_31260_1092# tinv7.ENB Do<5> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X31 a_36700_1090# a_35760_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X32 VDD a_35860_140# a_35760_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X33 VSS CLK cgate0.latch0.I1.ENB VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X34 a_14490_1090# Di<1> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X35 VDD a_15420_680# tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X36 a_16860_306# tinv7.EN Do<1> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X37 cgate0.nand0.OUT cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X38 dff_7.CLK cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X39 cgate0.latch0.I2.I CLK a_3720_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X40 a_25060_140# a_25390_140# a_25290_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X41 a_15210_190# a_14590_140# a_15100_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X42 VSS tinv0.I a_13260_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X43 a_29500_190# a_28560_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X44 a_10990_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X45 a_24060_306# tinv7.EN Do<3> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X46 VSS tinv7.I a_38460_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X47 a_33210_190# dff_7.CLK a_33100_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X48 VDD a_33420_680# a_33380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X49 dff_7.CLK cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X50 a_10990_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X51 cgate0.nand0.OUT cgate0.nand0.A a_5340_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X52 a_36190_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X53 cgate0.latch0.I1.ENB CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X54 a_11500_190# a_10560_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X55 a_32260_140# a_32590_140# a_32490_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X56 a_36190_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X57 a_26010_190# a_25390_140# a_25900_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X58 a_36700_190# a_35760_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X59 cgate0.latch0.I1.ENB CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X60 VSS cgate0.latch0.I2.I cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X61 a_21790_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X62 VSS tinv2.I a_20460_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X63 a_31260_306# tinv7.EN Do<5> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X64 dff_7.CLK cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X65 Do<1> tinv7.EN a_16860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X66 a_29780_1090# dff_7.CLK a_29610_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X67 VSS a_29820_680# a_29780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X68 tinv7.EN tinv7.ENB VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X69 a_22620_680# a_22410_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X70 a_32260_140# dff_7.CLK a_32490_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X71 a_11220_1090# a_10990_140# a_10660_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X72 VSS cgate0.nand0.OUT dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X73 a_3720_306# cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X74 a_15420_680# a_15210_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X75 Do<3> tinv7.ENB a_24060_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X76 a_36420_1090# a_36190_140# a_35860_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X77 nand.OUT WE a_300_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X78 a_36090_190# Di<7> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X79 tinv7.ENB RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X80 VSS a_11820_680# a_11780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X81 Do<3> tinv7.EN a_24060_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X82 a_33420_680# a_33210_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X83 a_27660_306# tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X84 a_22020_1090# a_21790_140# a_21460_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X85 VDD a_33420_680# tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X86 a_32490_1090# Di<6> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X87 VSS inv_and.O a_2460_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X88 a_13260_1092# tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X89 a_18420_190# dff_7.CLK a_17860_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X90 dff_7.O tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X91 VDD cgate0.nand0.OUT dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X92 VDD tinv4.I a_27660_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X93 VSS a_21360_190# a_22020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X94 dff_7.O tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X95 cgate0.nand0.A cgate0.latch0.I2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X96 a_34860_306# tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X97 a_38460_1092# tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X98 Do<5> tinv7.EN a_31260_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X99 VSS a_28660_140# a_28560_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X100 a_26180_190# a_25390_140# a_26010_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X101 VDD CLK cgate0.latch0.I1.ENB VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X102 dff_3.O tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X103 a_33210_190# a_32590_140# a_33100_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X104 VSS tinv7.ENB tinv7.EN VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X105 dff_2.O tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X106 a_28990_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X107 dff_7.CLK cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X108 a_25620_190# dff_7.CLK a_25060_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X109 VSS a_10660_140# a_10560_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X110 VDD a_24960_190# a_25620_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X111 VDD cgate0.nand0.OUT dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X112 VDD tinv7.ENB tinv7.EN VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X113 VSS a_35860_140# a_35760_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X114 a_33380_190# a_32590_140# a_33210_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X115 a_38460_1092# tinv7.ENB Do<7> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X116 VDD inv_and.O a_2460_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X117 a_300_306# SEL VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X118 VSS RE tinv7.ENB VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X119 a_22580_1090# dff_7.CLK a_22410_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X120 a_18810_190# dff_7.CLK a_18700_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X121 VSS CLK a_5340_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X122 VSS a_11820_680# tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X123 a_24060_1092# tinv7.ENB Do<3> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X124 a_29500_1090# a_28560_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X125 VDD a_28660_140# a_28560_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X126 VSS a_37020_680# tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X127 a_32820_190# dff_7.CLK a_32260_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X128 VDD RE tinv7.ENB VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X129 VSS cgate0.nand0.OUT dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X130 a_26010_190# dff_7.CLK a_25900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X131 VDD a_19020_680# tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X132 a_27660_306# tinv7.EN Do<4> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X133 dff_7.CLK cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X134 tinv7.EN tinv7.ENB VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X135 VDD tinv2.I a_20460_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X136 VDD a_26220_680# a_26180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X137 a_31260_1092# tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X138 a_35860_140# a_36190_140# a_36090_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X139 a_15100_190# a_14160_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X140 VDD a_11820_680# a_11780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X141 tinv7.ENB RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X142 VSS tinv7.ENB tinv7.EN VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X143 VSS tinv3.I a_24060_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X144 a_5340_306# CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X145 a_18810_190# a_18190_140# a_18700_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X146 a_34860_306# tinv7.EN Do<6> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X147 a_14590_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X148 dff_7.CLK cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X149 a_25060_140# dff_7.CLK a_25290_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X150 a_22300_190# a_21360_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X151 a_28890_190# Di<5> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X152 a_19020_680# a_18810_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X153 VSS tinv5.I a_31260_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X154 a_10660_140# dff_7.CLK a_10890_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X155 Do<1> tinv7.ENB a_16860_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X156 VSS a_15420_680# a_15380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X157 VDD a_21460_140# a_21360_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X158 a_22300_1090# a_21360_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X159 a_28990_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X160 tinv7.ENB RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X161 a_29220_1090# a_28990_140# a_28660_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X162 Do<4> tinv7.EN a_27660_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X163 a_26220_680# a_26010_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X164 a_14820_1090# a_14590_140# a_14260_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X165 a_10890_190# Di<0> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X166 VSS a_14160_190# a_14820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X167 a_25290_1090# Di<4> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X168 VDD a_26220_680# tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X169 a_18980_190# a_18190_140# a_18810_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X170 a_26220_680# a_26010_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X171 a_10890_1090# Di<0> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X172 tinv7.EN tinv7.ENB VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X173 a_13260_306# tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X174 a_38460_306# tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X175 inv_and.O nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X176 VDD a_11820_680# tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X177 VSS RE tinv7.ENB VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X178 dff_0.O tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X179 VSS a_22620_680# a_22580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X180 Do<6> tinv7.EN a_34860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X181 dff_1.O tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X182 VDD a_37020_680# tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X183 VSS cgate0.nand0.OUT dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X184 a_16860_1092# tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X185 a_33420_680# a_33210_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X186 a_29220_190# dff_7.CLK a_28660_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X187 a_11610_190# a_10990_140# a_11500_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X188 VSS a_14260_140# a_14160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X189 a_20460_306# tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X190 VDD a_17760_190# a_18420_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X191 cgate0.latch0.I2.I CLK a_2460_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X192 a_36810_190# a_36190_140# a_36700_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X193 a_15380_1090# dff_7.CLK a_15210_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X194 VSS a_15420_680# tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X195 a_16860_1092# tinv7.ENB Do<1> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X196 a_11220_190# dff_7.CLK a_10660_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X197 a_36420_190# dff_7.CLK a_35860_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X198 a_32590_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X199 VDD cgate0.nand0.A cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X200 VDD RE tinv7.ENB VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X201 VSS a_21460_140# a_21360_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X202 tinv7.EN tinv7.ENB VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X203 VDD nand.OUT inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X204 a_3720_1092# cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X205 a_29610_190# dff_7.CLK a_29500_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X206 a_2460_306# inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X207 VSS a_22620_680# tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X208 Do<6> tinv7.ENB a_34860_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X209 Do<2> tinv7.ENB a_20460_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X210 a_28660_140# a_28990_140# a_28890_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X211 VDD tinv0.I a_13260_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X212 a_11610_190# dff_7.CLK a_11500_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X213 VDD a_19020_680# a_18980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X214 VSS tinv1.I a_16860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X215 a_32820_1090# a_32590_140# a_32260_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X216 a_14590_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X217 a_36810_190# dff_7.CLK a_36700_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X218 a_24060_1092# tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X219 VDD tinv7.I a_38460_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X220 VSS a_29820_680# tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X221 a_10660_140# a_10990_140# a_10890_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X222 VDD a_29820_680# tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X223 a_38460_306# tinv7.EN Do<7> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X224 VDD a_29820_680# a_29780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X225 dff_6.O tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X226 VDD a_10560_190# a_11220_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X227 a_21790_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X228 a_34860_1092# tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X229 a_17860_140# dff_7.CLK a_18090_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X230 a_20460_306# tinv7.EN Do<2> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X231 VSS a_19020_680# a_18980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X232 VDD a_35760_190# a_36420_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X233 tinv7.ENB RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X234 VDD tinv7.ENB tinv7.EN VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X235 VDD a_14260_140# a_14160_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X236 a_15100_1090# a_14160_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X237 a_33380_1090# dff_7.CLK a_33210_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X238 cgate0.latch0.I2.I cgate0.latch0.I1.ENB a_3720_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X239 a_19020_680# a_18810_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X240 a_14490_190# Di<1> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X241 VSS a_17760_190# a_18420_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X242 a_28660_140# dff_7.CLK a_28890_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X243 a_33100_190# a_32160_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X244 a_34860_1092# tinv7.ENB Do<6> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X245 inv_and.O nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X246 VSS nand.OUT inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X247 a_18090_1090# Di<2> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X248 a_25900_1090# a_24960_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X249 VSS a_26220_680# a_26180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X250 tinv7.EN tinv7.ENB VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X251 dff_1.O tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X252 a_2460_306# cgate0.latch0.I1.ENB cgate0.latch0.I2.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X253 cgate0.nand0.A cgate0.latch0.I2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X254 a_11820_680# a_11610_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X255 a_21690_190# Di<3> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X256 a_28890_1090# Di<5> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X257 VSS a_24960_190# a_25620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X258 a_37020_680# a_36810_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X259 a_29780_190# a_28990_140# a_29610_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X260 a_24060_306# tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X261 VDD tinv5.I a_31260_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X262 VSS a_33420_680# a_33380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X263 VDD a_37020_680# a_36980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X264 dff_3.O tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X265 VDD a_22620_680# a_22580_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X266 cgate0.nand0.OUT CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X267 a_29610_190# a_28990_140# a_29500_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X268 VSS a_32160_190# a_32820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X269 a_11780_190# a_10990_140# a_11610_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X270 a_36980_190# a_36190_140# a_36810_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X271 VDD SEL nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X272 a_25390_140# dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X273 VSS a_25060_140# a_24960_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X274 a_31260_306# tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X275 dff_5.O tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X276 a_35860_140# dff_7.CLK a_36090_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X277 a_5340_306# cgate0.nand0.A cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X278 a_18980_1090# dff_7.CLK a_18810_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X279 a_33100_1090# a_32160_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X280 VSS a_26220_680# tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X281 a_11820_680# a_11610_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X282 a_21460_140# dff_7.CLK a_21690_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X283 Do<4> tinv7.ENB a_27660_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X284 VDD a_32260_140# a_32160_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X285 VDD tinv7.ENB tinv7.EN VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X286 tinv7.ENB RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X287 VSS a_32260_140# a_32160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X288 Do<0> tinv7.ENB a_13260_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X289 a_15210_190# dff_7.CLK a_15100_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X290 a_37020_680# a_36810_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X291 VDD cgate0.latch0.I2.I cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X292 a_18190_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X293 a_25620_1090# a_25390_140# a_25060_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X294 a_36090_1090# Di<7> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X295 VSS tinv7.ENB tinv7.EN VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X296 VSS a_33420_680# tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X297 Do<7> tinv7.ENB a_38460_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X298 a_14260_140# a_14590_140# a_14490_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X299 a_21690_1090# Di<3> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X300 VDD a_22620_680# tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X301 a_18700_190# a_17760_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X302 a_13260_306# tinv7.EN Do<0> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X303 a_22410_190# dff_7.CLK a_22300_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X304 VSS tinv4.I a_27660_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X305 VDD CLK cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X306 VSS RE tinv7.ENB VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X307 VDD tinv1.I a_16860_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X308 dff_4.O tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X309 a_25390_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X310 tinv7.ENB RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X311 a_27660_1092# tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X312 nand.OUT WE VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X313 a_22410_190# a_21790_140# a_22300_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X314 a_21460_140# a_21790_140# a_21690_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X315 dff_0.O tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X316 VDD a_28560_190# a_29220_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X317 a_25900_190# a_24960_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X318 a_18090_190# Di<2> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X319 VSS tinv6.I a_34860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X320 a_26180_1090# dff_7.CLK a_26010_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X321 a_32590_140# dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X322 VDD a_14160_190# a_14820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X323 a_27660_1092# tinv7.ENB Do<4> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X324 a_11780_1090# dff_7.CLK a_11610_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X325 tinv7.EN tinv7.ENB VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X326 a_18700_1090# a_17760_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X327 a_2460_1092# inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X328 a_13260_1092# tinv7.ENB Do<0> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X329 VDD a_17860_140# a_17760_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X330 a_29820_680# a_29610_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X331 a_25290_190# Di<4> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X332 a_36980_1090# dff_7.CLK a_36810_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X333 Do<0> tinv7.EN a_13260_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X334 a_16860_306# tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X335 VSS a_28560_190# a_29220_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X336 Do<7> tinv7.EN a_38460_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X337 Do<5> tinv7.ENB a_31260_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X338 VSS a_37020_680# a_36980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X339 VDD tinv3.I a_24060_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X340 dff_4.O tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X341 a_2460_1092# CLK cgate0.latch0.I2.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X342 VSS a_10560_190# a_11220_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X343 a_32490_190# Di<6> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
.ends

