magic
tech gf180mcuC
magscale 1 10
timestamp 1684461354
<< nwell >>
rect -150 -90 330 570
<< pmos >>
rect 60 136 120 476
<< pdiff >>
rect -60 450 60 476
rect -60 390 -31 450
rect 31 390 60 450
rect -60 330 60 390
rect -60 270 -31 330
rect 31 270 60 330
rect -60 210 60 270
rect -60 150 -31 210
rect 31 150 60 210
rect -60 136 60 150
rect 120 450 240 476
rect 120 390 149 450
rect 211 390 240 450
rect 120 330 240 390
rect 120 270 149 330
rect 211 270 240 330
rect 120 210 240 270
rect 120 150 149 210
rect 211 150 240 210
rect 120 136 240 150
<< pdiffc >>
rect -31 390 31 450
rect -31 270 31 330
rect -31 150 31 210
rect 149 390 211 450
rect 149 270 211 330
rect 149 150 211 210
<< polysilicon >>
rect 4 650 120 666
rect 4 580 20 650
rect 70 580 120 650
rect 4 564 120 580
rect 60 476 120 564
rect 60 84 120 136
<< polycontact >>
rect 20 580 70 650
<< metal1 >>
rect -44 650 86 672
rect -44 580 20 650
rect 70 580 86 650
rect -44 560 86 580
rect -44 450 44 476
rect -44 390 -31 450
rect 31 390 44 450
rect -44 330 44 390
rect -44 270 -31 330
rect 31 270 44 330
rect -44 210 44 270
rect -44 150 -31 210
rect 31 150 44 210
rect -44 136 44 150
rect 136 450 224 476
rect 136 390 149 450
rect 211 390 224 450
rect 136 330 224 390
rect 136 270 149 330
rect 211 270 224 330
rect 136 210 224 270
rect 136 150 149 210
rect 211 150 224 210
rect 136 136 224 150
<< end >>
