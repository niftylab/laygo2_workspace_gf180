magic
tech gf180mcuC
magscale 1 10
timestamp 1683427464
<< nmos >>
rect 60 306 120 476
<< ndiff >>
rect -60 459 60 476
rect -60 413 -30 459
rect 30 413 60 459
rect -60 365 60 413
rect -60 319 -30 365
rect 30 319 60 365
rect -60 306 60 319
rect 120 459 240 476
rect 120 413 150 459
rect 210 413 240 459
rect 120 365 240 413
rect 120 319 150 365
rect 210 319 240 365
rect 120 306 240 319
<< ndiffc >>
rect -30 413 30 459
rect -30 319 30 365
rect 150 413 210 459
rect 150 319 210 365
<< polysilicon >>
rect -44 650 120 666
rect -44 580 -30 650
rect 30 580 120 650
rect -44 566 120 580
rect 60 476 120 566
rect 60 262 120 306
<< polycontact >>
rect -30 580 30 650
<< metal1 >>
rect -44 650 44 672
rect -44 580 -30 650
rect 30 580 44 650
rect -44 560 44 580
rect -44 459 44 476
rect -44 413 -30 459
rect 30 413 44 459
rect -44 365 44 413
rect -44 319 -30 365
rect 30 319 44 365
rect -44 280 44 319
rect 136 459 224 476
rect 136 413 150 459
rect 210 413 224 459
rect 136 365 224 413
rect 136 319 150 365
rect 210 319 224 365
rect 136 280 224 319
<< end >>
