* NGSPICE file created from dff_byte_left.ext - technology: gf180mcuC

.subckt dff_byte_left CLK Di<0> Di<1> Di<2> Di<3> Di<4> Di<5> Di<6> Di<7> Do<0> Do<1>
+ Do<2> Do<3> Do<4> Do<5> Do<6> Do<7> RE SEL WE VSS VDD
X0 a_1380_680# a_1170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1 VSS a_1380_680# tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2 a_19380_680# a_19170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3 VSS tinv5.I a_20820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4 VSS CLK cgate0.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5 a_7980_1090# a_7750_140# a_7420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6 a_7420_140# a_7750_140# a_7650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7 a_11020_140# cgate0.inv1.O a_11250_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8 VSS a_15780_680# a_15740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9 Do<4> buf_RE1.O a_17220_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10 VDD cgate0.latch0.I2.I cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11 cgate0.inv1.O cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12 a_15740_1090# cgate0.inv1.O a_15570_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X13 VDD a_4980_680# tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X14 a_15180_1090# a_14950_140# a_14620_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X15 a_17220_1092# buf_RE0.O Do<4> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X16 a_6420_1092# tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X17 a_4150_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X18 Do<7> buf_RE0.O a_28020_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X19 a_13620_306# tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X20 VSS a_14520_190# a_15180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X21 VDD a_12180_680# tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X22 Do<6> buf_RE1.O a_24420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X23 VSS a_22980_680# a_22940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X24 a_4770_190# a_4150_140# a_4660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X25 VSS tinv0.I a_2820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X26 a_25980_1090# a_25750_140# a_25420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X27 a_6420_1092# buf_RE0.O Do<1> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X28 a_18780_190# cgate0.inv1.O a_18220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X29 a_220_140# cgate0.inv1.O a_450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X30 VDD a_19380_680# a_19340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X31 VDD a_22980_680# tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X32 a_20820_306# tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X33 buf_RE1.O buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X34 cgate0.inv0.O CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X35 VSS a_21720_190# a_22380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X36 a_12140_190# a_11350_140# a_11970_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X37 a_24420_1092# tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X38 Do<0> buf_RE0.O a_2820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X39 VSS a_4980_680# a_4940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X40 Do<1> buf_RE1.O a_6420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X41 a_25980_190# cgate0.inv1.O a_25420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X42 a_22770_190# a_22150_140# a_22660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X43 VDD buf_RE0.O buf_RE1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X44 VDD cgate0.nand0.OUT cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X45 a_780_190# cgate0.inv1.O a_220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X46 a_24420_1092# buf_RE0.O Do<6> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X47 VSS nand.OUT inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X48 VDD tinv1.I a_6420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X49 a_2820_306# tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X50 VSS a_3720_190# a_4380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X51 a_10020_1092# buf_RE0.O Do<2> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X52 Do<5> buf_RE0.O a_20820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X53 a_19380_680# a_19170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X54 VDD cgate0.nand0.A a_35760_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X55 a_7980_190# cgate0.inv1.O a_7420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X56 a_18450_1090# Di<5> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X57 VDD a_4980_680# a_4940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X58 a_14950_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X59 VSS tinv4.I a_17220_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X60 VDD a_3720_190# a_4380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X61 a_1340_190# a_550_140# a_1170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X62 a_13620_306# buf_RE1.O Do<3> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X63 VDD buf_RE0.O buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X64 a_7750_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X65 cgate0.nand0.OUT CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X66 a_8260_1090# a_7320_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X67 VDD a_12180_680# a_12140_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X68 a_11020_140# a_11350_140# a_11250_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X69 VDD tinv6.I a_24420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X70 VSS RE buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X71 VDD a_7420_140# a_7320_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X72 a_8580_680# a_8370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X73 a_15460_190# a_14520_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X74 VSS tinv6.I a_24420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X75 a_20820_306# buf_RE1.O Do<5> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X76 cgate0.inv1.O cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X77 VDD a_22980_680# a_22940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X78 VSS a_19380_680# a_19340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X79 cgate0.inv1.O cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X80 a_14850_190# Di<4> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X81 VDD a_21720_190# a_22380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X82 a_22660_190# a_21720_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X83 a_25750_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X84 cgate0.nand0.A cgate0.latch0.I2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X85 inv_and.O nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X86 a_4050_1090# Di<1> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X87 a_17220_306# tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X88 a_26260_1090# a_25320_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X89 a_26580_680# a_26370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X90 buf_RE0.O RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X91 a_14620_140# cgate0.inv1.O a_14850_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X92 dff_4.O tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X93 VDD a_25420_140# a_25320_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X94 Do<7> buf_RE1.O a_28020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X95 VSS a_26580_680# a_26540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X96 cgate0.nand0.OUT cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X97 a_1170_190# cgate0.inv1.O a_1060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X98 VSS tinv1.I a_6420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X99 a_33420_306# cgate0.nand0.A cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X100 a_2820_306# buf_RE1.O Do<0> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X101 dff_2.O tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X102 a_11860_1090# a_10920_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X103 a_12180_680# a_11970_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X104 a_12180_680# a_11970_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X105 buf_RE0.O RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X106 a_22050_190# Di<6> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X107 a_10020_1092# tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X108 a_11250_1090# Di<3> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X109 a_18780_1090# a_18550_140# a_18220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X110 VDD WE nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X111 Do<2> buf_RE1.O a_10020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X112 VSS a_25320_190# a_25980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X113 a_24420_306# tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X114 a_4660_190# a_3720_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X115 a_35760_306# CLK cgate0.latch0.I2.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X116 VSS cgate0.nand0.OUT cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X117 VDD CLK cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X118 a_550_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X119 a_3820_140# cgate0.inv1.O a_4050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X120 VDD a_15780_680# tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X121 dff_6.O tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X122 a_1060_1090# a_120_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X123 a_8540_1090# cgate0.inv1.O a_8370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X124 a_17220_1092# tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X125 a_22050_1090# Di<6> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X126 VSS buf_RE0.O buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X127 VSS a_8580_680# a_8540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X128 VSS a_14620_140# a_14520_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X129 VSS RE buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X130 a_4050_190# Di<1> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X131 a_15570_190# a_14950_140# a_15460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X132 dff_7.O tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X133 a_28020_1092# tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X134 a_450_1090# Di<0> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X135 Do<1> buf_RE0.O a_6420_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X136 a_6420_306# tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X137 VSS a_7320_190# a_7980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X138 a_11580_190# cgate0.inv1.O a_11020_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X139 VSS a_15780_680# tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X140 a_36300_306# cgate0.inv0.O cgate0.latch0.I2.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X141 dff_1.O tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X142 a_21820_140# cgate0.inv1.O a_22050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X143 VDD RE buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X144 cgate0.nand0.OUT cgate0.nand0.A a_33420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X145 VSS a_21820_140# a_21720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X146 VDD cgate0.nand0.A cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X147 a_1380_680# a_1170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X148 Do<3> buf_RE0.O a_13620_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X149 a_26540_1090# cgate0.inv1.O a_26370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X150 a_28020_1092# buf_RE0.O Do<7> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X151 cgate0.inv1.O cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X152 a_18550_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X153 VSS a_22980_680# tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X154 nand.OUT SEL VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X155 dff_0.O tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X156 a_11580_1090# a_11350_140# a_11020_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X157 buf_RE1.O buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X158 a_2820_1092# tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X159 a_11970_190# cgate0.inv1.O a_11860_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X160 Do<6> buf_RE0.O a_24420_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X161 a_19060_190# a_18120_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X162 buf_RE0.O RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X163 a_36300_1092# inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X164 VDD tinv4.I a_17220_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X165 a_1340_1090# cgate0.inv1.O a_1170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X166 VSS a_3820_140# a_3720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X167 VSS tinv7.I a_28020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X168 a_25750_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X169 cgate0.latch0.I2.I cgate0.inv0.O a_36300_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X170 a_24420_306# buf_RE1.O Do<6> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X171 a_2820_1092# buf_RE0.O Do<0> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X172 VSS a_4980_680# tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X173 VDD a_15780_680# a_15740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X174 a_21820_140# a_22150_140# a_22050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X175 cgate0.inv0.O CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X176 VSS tinv2.I a_10020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X177 dff_5.O tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X178 a_18450_190# Di<5> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X179 inv_and.O nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X180 a_26260_190# a_25320_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X181 a_780_1090# a_550_140# a_220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X182 VDD a_14520_190# a_15180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X183 a_20820_1092# tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X184 a_18550_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X185 VSS cgate0.nand0.OUT cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X186 a_19060_1090# a_18120_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X187 a_6420_306# buf_RE1.O Do<1> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X188 a_7750_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X189 VDD a_18220_140# a_18120_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X190 a_15780_680# a_15570_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X191 VSS a_18120_190# a_18780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X192 VSS CLK a_33420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X193 a_25650_190# Di<7> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X194 a_3820_140# a_4150_140# a_4050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X195 a_20820_1092# buf_RE0.O Do<5> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X196 VDD tinv0.I a_2820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X197 VSS a_12180_680# a_12140_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X198 Do<3> buf_RE1.O a_13620_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X199 cgate0.inv1.O cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X200 a_450_190# Di<0> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X201 a_8260_190# a_7320_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X202 VSS SEL a_39180_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X203 dff_7.O tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X204 buf_RE1.O buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X205 a_22980_680# a_22770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X206 VDD tinv2.I a_10020_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X207 a_14850_1090# Di<4> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X208 a_15740_190# a_14950_140# a_15570_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X209 VSS a_18220_140# a_18120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X210 Do<5> buf_RE1.O a_20820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X211 VSS a_120_190# a_780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X212 a_7650_190# Di<2> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X213 VDD CLK cgate0.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X214 a_7420_140# cgate0.inv1.O a_7650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X215 a_4660_1090# a_3720_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X216 VDD tinv5.I a_20820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X217 a_15180_190# cgate0.inv1.O a_14620_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X218 VSS inv_and.O a_36300_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X219 VDD a_3820_140# a_3720_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X220 a_4980_680# a_4770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X221 dff_2.O tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X222 a_33420_306# CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X223 a_22940_190# a_22150_140# a_22770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X224 VSS a_25420_140# a_25320_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X225 a_4980_680# a_4770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X226 a_11350_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X227 VDD nand.OUT inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X228 VDD a_8580_680# tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X229 a_19340_1090# cgate0.inv1.O a_19170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X230 a_39180_306# WE nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X231 VSS a_220_140# a_120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X232 VSS a_1380_680# a_1340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X233 Do<0> buf_RE1.O a_2820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X234 VDD a_11020_140# a_10920_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X235 VSS a_26580_680# tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X236 a_22380_190# cgate0.inv1.O a_21820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X237 a_25420_140# cgate0.inv1.O a_25650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X238 cgate0.nand0.A cgate0.latch0.I2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X239 a_15570_190# cgate0.inv1.O a_15460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X240 a_22660_1090# a_21720_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X241 a_22980_680# a_22770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X242 a_8370_190# a_7750_140# a_8260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X243 a_4940_190# a_4150_140# a_4770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X244 Do<4> buf_RE0.O a_17220_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X245 a_17220_306# buf_RE1.O Do<4> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X246 VDD a_21820_140# a_21720_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X247 VDD buf_RE0.O buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X248 VSS a_7420_140# a_7320_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X249 dff_1.O tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X250 a_14620_140# a_14950_140# a_14850_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X251 VDD cgate0.nand0.OUT cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X252 VDD a_26580_680# tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X253 a_4380_190# cgate0.inv1.O a_3820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X254 VSS a_8580_680# tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X255 a_22770_190# cgate0.inv1.O a_22660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X256 VDD a_220_140# a_120_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X257 a_11350_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X258 buf_RE0.O RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X259 dff_3.O tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X260 a_4940_1090# cgate0.inv1.O a_4770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X261 a_13620_1092# tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X262 a_4380_1090# a_4150_140# a_3820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X263 a_26370_190# a_25750_140# a_26260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X264 a_11970_190# a_11350_140# a_11860_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X265 a_12140_1090# cgate0.inv1.O a_11970_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X266 dff_6.O tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X267 buf_RE0.O RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X268 VDD a_1380_680# tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X269 VDD a_18120_190# a_18780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X270 a_4770_190# cgate0.inv1.O a_4660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X271 a_13620_1092# buf_RE0.O Do<3> VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X272 a_11250_190# Di<3> VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X273 buf_RE1.O buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X274 VDD a_8580_680# a_8540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X275 Do<2> buf_RE0.O a_10020_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X276 a_22940_1090# cgate0.inv1.O a_22770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X277 VSS RE buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X278 a_28020_306# tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X279 a_26580_680# a_26370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X280 a_1170_190# a_550_140# a_1060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X281 a_22380_1090# a_22150_140# a_21820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X282 a_19340_190# a_18550_140# a_19170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X283 VDD a_7320_190# a_7980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X284 a_35760_1092# cgate0.inv0.O cgate0.latch0.I2.I VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X285 a_550_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X286 dff_3.O tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X287 buf_RE1.O buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X288 VSS a_10920_190# a_11580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X289 VDD a_19380_680# tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X290 VDD tinv7.I a_28020_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X291 VDD RE buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X292 VSS buf_RE0.O buf_RE1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X293 VDD tinv3.I a_13620_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X294 a_26540_190# a_25750_140# a_26370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X295 a_1060_190# a_120_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X296 cgate0.inv1.O cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X297 cgate0.latch0.I2.I CLK a_36300_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X298 a_8580_680# a_8370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X299 a_10020_306# tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X300 dff_5.O tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X301 VDD a_26580_680# a_26540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X302 VDD a_25320_190# a_25980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X303 VDD RE buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X304 VSS a_11020_140# a_10920_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X305 buf_RE0.O RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X306 a_7650_1090# Di<2> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X307 VDD a_10920_190# a_11580_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X308 a_19170_190# cgate0.inv1.O a_19060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X309 VDD inv_and.O a_36300_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X310 a_14950_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X311 a_18220_140# cgate0.inv1.O a_18450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X312 a_8540_190# a_7750_140# a_8370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X313 a_15460_1090# a_14520_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X314 VSS a_12180_680# tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X315 VSS cgate0.nand0.OUT cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X316 VDD cgate0.nand0.OUT cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X317 VDD a_14620_140# a_14520_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X318 a_15780_680# a_15570_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X319 a_18220_140# a_18550_140# a_18450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X320 VSS buf_RE0.O buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X321 VDD a_1380_680# a_1340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X322 dff_0.O tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X323 VSS cgate0.latch0.I2.I cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X324 a_28020_306# buf_RE1.O Do<7> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X325 a_26370_190# cgate0.inv1.O a_26260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X326 a_4150_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X327 VSS a_19380_680# tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X328 a_25650_1090# Di<7> VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X329 a_36300_306# inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X330 a_25420_140# a_25750_140# a_25650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X331 VDD a_120_190# a_780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X332 VSS tinv3.I a_13620_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X333 a_36300_1092# CLK cgate0.latch0.I2.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X334 a_10020_306# buf_RE1.O Do<2> VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X335 a_19170_190# a_18550_140# a_19060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X336 VSS cgate0.nand0.A a_35760_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X337 a_220_140# a_550_140# a_450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X338 a_22150_140# cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X339 a_8370_190# cgate0.inv1.O a_8260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X340 dff_4.O tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X341 a_11860_190# a_10920_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X342 a_22150_140# cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X343 buf_RE1.O buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
.ends

