** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/RAM8.sch
.subckt RAM8 Di0 Do0_buf Di1 Do1_buf Di2 Do2_buf Di3 Do3_buf Di4 Do4_buf Di5 Do5_buf Di6 Do6_buf Di7
+ Do7_buf Di8 Do8_buf Di9 Do9_buf Di10 Do10_buf Di11 Do11_buf Di12 Do12_buf Di13 Do13_buf Di14 Do14_buf Di15
+ Do15_buf Di16 Do16_buf Di17 Do17_buf Di18 Do18_buf Di19 Do19_buf Di20 Do20_buf Di21 Do21_buf Di22 Do22_buf
+ Di23 Do23_buf Di24 Do24_buf Di25 Do25_buf Di26 Do26_buf Di27 Do27_buf Di28 Do28_buf Di29 Do29_buf Di30
+ Do30_buf Di31 Do31_buf VDD VSS WE0 WE1 WE2 WE3 CLK A0 A1 A2 EN RE
*.PININFO Di0:I Do0_buf:O Di1:I Do1_buf:O Di2:I Do2_buf:O Di3:I Do3_buf:O Di4:I Do4_buf:O Di5:I
*+ Do5_buf:O Di6:I Do6_buf:O Di7:I Do7_buf:O Di8:I Do8_buf:O Di9:I Do9_buf:O Di10:I Do10_buf:O Di11:I Do11_buf:O
*+ Di12:I Do12_buf:O Di13:I Do13_buf:O Di14:I Do14_buf:O Di15:I Do15_buf:O Di16:I Do16_buf:O Di17:I
*+ Do17_buf:O Di18:I Do18_buf:O Di19:I Do19_buf:O Di20:I Do20_buf:O Di21:I Do21_buf:O Di22:I Do22_buf:O Di23:I
*+ Do23_buf:O Di24:I Do24_buf:O Di25:I Do25_buf:O Di26:I Do26_buf:O Di27:I Do27_buf:O Di28:I Do28_buf:O Di29:I
*+ Do29_buf:O Di30:I Do30_buf:O Di31:I Do31_buf:O VDD:B VSS:B WE0:I WE1:I WE2:I WE3:I CLK:I A0:I A1:I A2:I EN:I
*+ RE:I
xbyte1 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL0 CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte2 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL1 CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte3 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL2 CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte4 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL[3] CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte5 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL[4] CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte6 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL[5] CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte7 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL[6] CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
xbyte8 VDD VSS we3_buf we2_buf we1_buf we0_buf SEL[7] CLK_buf di9_buf di7_buf Di[19] Di[20] Di[30]
+ di8_buf di10_buf di4_buf di12_buf Di[24] di5_buf Di[23] Di[29] di3_buf di14_buf Di[18] Di[28] Di[17]
+ di16_buf Di[27] Di[21] Di[22] di0_buf di1_buf Di[31] Di[26] Di[25] di15_buf di2_buf di13_buf di6_buf
+ di11_buf Do21 Do22 Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6
+ Do5 Do18 Do0 Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE_buf word NF=2
x_dec1 A1 EN A2 A0 VDD VSS Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 dec_3to8 NF=2
X_inv1 Y0 VDD VSS net1 inv NF=2
X_inv2 net1 VDD VSS SEL0 inv NF=8
X_inv3 Y1 VDD VSS net2 inv NF=2
X_inv4 net2 VDD VSS SEL1 inv NF=8
X_inv65 net9 VDD VSS CLK_buf inv NF=8
X_inv73 WE0 VDD VSS net13 inv NF=1
X_inv74 net13 VDD VSS we0_buf inv NF=4
X_inv75 Di0 VDD VSS net14 inv NF=2
X_inv76 net14 VDD VSS di0_buf inv NF=8
X_inv143 CLK VDD VSS net9 inv NF=2
X_inv9 Y4 VDD VSS net5 inv NF=2
X_inv10 net5 VDD VSS SEL[4] inv NF=8
X_inv11 Y5 VDD VSS net6 inv NF=2
X_inv36 net6 VDD VSS SEL[5] inv NF=8
X_inv5 Y2 VDD VSS net3 inv NF=2
X_inv13 Y6 VDD VSS net7 inv NF=2
X_inv6 net3 VDD VSS SEL2 inv NF=8
X_inv14 net7 VDD VSS SEL[6] inv NF=8
X_inv7 Y3 VDD VSS net4 inv NF=2
X_inv15 Y7 VDD VSS net8 inv NF=2
X_inv8 net4 VDD VSS SEL[3] inv NF=8
X_inv16 net8 VDD VSS SEL[7] inv NF=8
X_inv67 WE1 VDD VSS net12 inv NF=1
X_inv68 WE2 VDD VSS net11 inv NF=1
X_inv69 WE3 VDD VSS net10 inv NF=1
X_inv70 net12 VDD VSS we1_buf inv NF=4
X_inv71 net11 VDD VSS we2_buf inv NF=4
X_inv72 net10 VDD VSS we3_buf inv NF=4
X_inv12 Do0 VDD VSS net46 inv NF=1
X_inv17 net46 VDD VSS Do0_buf inv NF=4
X_inv32 Do8 VDD VSS net47 inv NF=1
X_inv33 net47 VDD VSS Do8_buf inv NF=4
X_inv49 Do16 VDD VSS net48 inv NF=1
X_inv50 net48 VDD VSS Do16_buf inv NF=4
X_inv66 Do24 VDD VSS net49 inv NF=1
X_inv139 net49 VDD VSS Do24_buf inv NF=4
X_inv18 Do1 VDD VSS net50 inv NF=1
X_inv19 net50 VDD VSS Do1_buf inv NF=4
X_inv20 Do2 VDD VSS net51 inv NF=1
X_inv21 net51 VDD VSS Do2_buf inv NF=4
X_inv22 Do3 VDD VSS net52 inv NF=1
X_inv23 net52 VDD VSS Do3_buf inv NF=4
X_inv24 Do4 VDD VSS net53 inv NF=1
X_inv25 net53 VDD VSS Do4_buf inv NF=4
X_inv26 Do5 VDD VSS net54 inv NF=1
X_inv27 net54 VDD VSS Do5_buf inv NF=4
X_inv28 Do6 VDD VSS net55 inv NF=1
X_inv29 net55 VDD VSS Do6_buf inv NF=4
X_inv30 Do7 VDD VSS net56 inv NF=1
X_inv31 net56 VDD VSS Do7_buf inv NF=4
X_inv34 Do9 VDD VSS net57 inv NF=1
X_inv35 net57 VDD VSS Do9_buf inv NF=4
X_inv37 Do10 VDD VSS net58 inv NF=1
X_inv38 net58 VDD VSS Do10_buf inv NF=4
X_inv39 Do11 VDD VSS net59 inv NF=1
X_inv40 net59 VDD VSS Do11_buf inv NF=4
X_inv41 Do12 VDD VSS net60 inv NF=1
X_inv42 net60 VDD VSS Do12_buf inv NF=4
X_inv43 Do13 VDD VSS net61 inv NF=1
X_inv44 net61 VDD VSS Do13_buf inv NF=4
X_inv45 Do14 VDD VSS net62 inv NF=1
X_inv46 net62 VDD VSS Do14_buf inv NF=4
X_inv47 Do15 VDD VSS net63 inv NF=1
X_inv48 net63 VDD VSS Do15_buf inv NF=4
X_inv51 Do17 VDD VSS net64 inv NF=1
X_inv52 net64 VDD VSS Do17_buf inv NF=4
X_inv53 Do18 VDD VSS net65 inv NF=1
X_inv54 net65 VDD VSS Do18_buf inv NF=4
X_inv55 Do19 VDD VSS net66 inv NF=1
X_inv56 net66 VDD VSS Do19_buf inv NF=4
X_inv57 Do20 VDD VSS net67 inv NF=1
X_inv58 net67 VDD VSS Do20_buf inv NF=4
X_inv59 Do21 VDD VSS net68 inv NF=1
X_inv60 net68 VDD VSS Do21_buf inv NF=4
X_inv61 Do22 VDD VSS net69 inv NF=1
X_inv62 net69 VDD VSS Do22_buf inv NF=4
X_inv63 Do23 VDD VSS net70 inv NF=1
X_inv64 net70 VDD VSS Do23_buf inv NF=4
X_inv140 Do25 VDD VSS net71 inv NF=1
X_inv141 net71 VDD VSS Do25_buf inv NF=4
X_inv142 Do26 VDD VSS net72 inv NF=1
X_inv144 net72 VDD VSS Do26_buf inv NF=4
X_inv145 Do27 VDD VSS net73 inv NF=1
X_inv146 net73 VDD VSS Do27_buf inv NF=4
X_inv147 Do28 VDD VSS net74 inv NF=1
X_inv148 net74 VDD VSS Do28_buf inv NF=4
X_inv149 Do29 VDD VSS net75 inv NF=1
X_inv150 net75 VDD VSS Do29_buf inv NF=4
X_inv151 Do30 VDD VSS net76 inv NF=1
X_inv152 net76 VDD VSS Do30_buf inv NF=4
X_inv153 Do31 VDD VSS net77 inv NF=1
X_inv154 net77 VDD VSS Do31_buf inv NF=4
X_inv83 Di4 VDD VSS net15 inv NF=2
X_inv91 Di8 VDD VSS net16 inv NF=2
X_inv99 Di12 VDD VSS net17 inv NF=2
X_inv115 Di16 VDD VSS net18 inv NF=2
X_inv107 Di20 VDD VSS net19 inv NF=2
X_inv123 Di24 VDD VSS net20 inv NF=2
X_inv131 Di28 VDD VSS net21 inv NF=2
X_inv77 Di1 VDD VSS net22 inv NF=2
X_inv85 Di5 VDD VSS net23 inv NF=2
X_inv86 Di9 VDD VSS net24 inv NF=2
X_inv93 Di13 VDD VSS net25 inv NF=2
X_inv94 Di17 VDD VSS net26 inv NF=2
X_inv101 Di21 VDD VSS net27 inv NF=2
X_inv102 Di25 VDD VSS net28 inv NF=2
X_inv109 Di29 VDD VSS net29 inv NF=2
X_inv84 net15 VDD VSS di4_buf inv NF=8
X_inv92 net16 VDD VSS di8_buf inv NF=8
X_inv100 net17 VDD VSS di12_buf inv NF=8
X_inv108 net18 VDD VSS di16_buf inv NF=8
X_inv116 net19 VDD VSS Di[20] inv NF=8
X_inv124 net20 VDD VSS Di[24] inv NF=8
X_inv132 net21 VDD VSS Di[28] inv NF=8
X_inv78 net22 VDD VSS di1_buf inv NF=8
X_inv110 net23 VDD VSS di5_buf inv NF=8
X_inv117 net24 VDD VSS di9_buf inv NF=8
X_inv118 net25 VDD VSS di13_buf inv NF=8
X_inv125 net26 VDD VSS Di[17] inv NF=8
X_inv126 net27 VDD VSS Di[21] inv NF=8
X_inv133 net28 VDD VSS Di[25] inv NF=8
X_inv134 net29 VDD VSS Di[29] inv NF=8
X_inv80 net30 VDD VSS di2_buf inv NF=8
X_inv96 net31 VDD VSS di6_buf inv NF=8
X_inv97 net32 VDD VSS di10_buf inv NF=8
X_inv98 net33 VDD VSS di14_buf inv NF=8
X_inv103 net34 VDD VSS Di[18] inv NF=8
X_inv104 net35 VDD VSS Di[22] inv NF=8
X_inv105 net36 VDD VSS Di[26] inv NF=8
X_inv106 net37 VDD VSS Di[30] inv NF=8
X_inv112 net38 VDD VSS di3_buf inv NF=8
X_inv128 net39 VDD VSS di7_buf inv NF=8
X_inv129 net40 VDD VSS di11_buf inv NF=8
X_inv130 net41 VDD VSS di15_buf inv NF=8
X_inv135 net42 VDD VSS Di[19] inv NF=8
X_inv136 net43 VDD VSS Di[23] inv NF=8
X_inv137 net44 VDD VSS Di[27] inv NF=8
X_inv138 net45 VDD VSS Di[31] inv NF=8
X_inv79 Di2 VDD VSS net30 inv NF=2
X_inv81 Di6 VDD VSS net31 inv NF=2
X_inv82 Di10 VDD VSS net32 inv NF=2
X_inv87 Di14 VDD VSS net33 inv NF=2
X_inv88 Di18 VDD VSS net34 inv NF=2
X_inv89 Di22 VDD VSS net35 inv NF=2
X_inv90 Di26 VDD VSS net36 inv NF=2
X_inv95 Di30 VDD VSS net37 inv NF=2
X_inv111 Di3 VDD VSS net38 inv NF=2
X_inv113 Di7 VDD VSS net39 inv NF=2
X_inv114 Di11 VDD VSS net40 inv NF=2
X_inv119 Di15 VDD VSS net41 inv NF=2
X_inv120 Di19 VDD VSS net42 inv NF=2
X_inv121 Di23 VDD VSS net43 inv NF=2
X_inv122 Di27 VDD VSS net44 inv NF=2
X_inv127 Di31 VDD VSS net45 inv NF=2
X_inv155 RE VDD VSS net78 inv NF=2
X_inv156 net78 VDD VSS RE_buf inv NF=8
.ends

* expanding   symbol:  xschem_lib/DFFRAM_full_custom/word.sym # of pins=73
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/word.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/word.sch
.subckt word  VDD VSS WE3 WE2 WE1 WE0 SEL CLK Di9 Di7 Di19 Di20 Di30 Di8 Di10 Di4 Di12 Di24 Di5 Di23
+ Di29 Di3 Di14 Di18 Di28 Di17 Di16 Di27 Di21 Di22 Di0 Di1 Di31 Di26 Di25 Di15 Di2 Di13 Di6 Di11 Do21 Do22
+ Do27 Do23 Do28 Do8 Do9 Do10 Do11 Do12 Do29 Do30 Do13 Do14 Do15 Do16 Do24 Do17 Do1 Do7 Do6 Do5 Do18 Do0
+ Do2 Do3 Do4 Do19 Do20 Do25 Do26 Do31 RE   NF=2
*.PININFO SEL:I WE0:I Di31:I Di30:I Di29:I Di28:I Di27:I Di26:I Di25:I Di24:I Do31:O Do30:O Do29:O
*+ Do28:O Do27:O Do26:O Do25:O Do24:O VDD:B VSS:B Di23:I Di22:I Di21:I Di20:I Di19:I Di18:I Di17:I Di16:I
*+ Do23:O Do22:O Do21:O Do20:O Do19:O Do18:O Do17:O Do16:O Di15:I Di14:I Di13:I Di12:I Di11:I Di10:I Di9:I
*+ Di8:I Do15:O Do14:O Do13:O Do12:O Do11:O Do10:O Do9:O Do8:O Di7:I Di6:I Di5:I Di4:I Di3:I Di2:I Di1:I
*+ Di0:I Do7:O Do6:O Do5:O Do4:O Do3:O Do2:O Do1:O Do0:O WE1:I WE2:I WE3:I CLK:I RE:I
xByte_1 VDD VSS WE0 Di3 Di7 Do3 Do7 CLK_buf SEL_buf Di2 Di6 Do2 Do6 Di5 Di1 Do5 Do1 Di4 Do4 Di0 Do0
+ RE_buf byte_dff NF=NF
X_inv1 SEL VDD VSS SEL_bar inv NF=1
X_inv2 SEL_bar VDD VSS SEL_buf inv NF=4
xByte_2 VDD VSS WE1 Di11 Di15 Do11 Do15 CLK_buf SEL_buf Di10 Di14 Do10 Do14 Di13 Di9 Do13 Do9 Di12
+ Do12 Di8 Do8 RE_buf byte_dff NF=NF
xByte_3 VDD VSS WE2 Di19 Di23 Do19 Do23 CLK_buf SEL_buf Di18 Di22 Do18 Do22 Di21 Di17 Do21 Do17 Di20
+ Do20 Di16 Do16 RE_buf byte_dff NF=NF
xByte_4 VDD VSS WE3 Di27 Di31 Do27 Do31 CLK_buf SEL_buf Di26 Di30 Do26 Do30 Di29 Di25 Do29 Do25 Di28
+ Do28 Di24 Do24 RE_buf byte_dff NF=NF
X_inv3 CLK VDD VSS CLK_bar inv NF=2
X_inv4 CLK_bar VDD VSS CLK_buf inv NF=8
X_inv5 net1 VDD VSS RE_bar inv NF=NF*3
X_inv6 RE_bar VDD VSS RE_buf inv NF=NF*9
X_nand1 RE SEL net2 VDD VSS nand NF=1
X_inv7 net2 VDD VSS net1 inv NF=NF
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/dec_3to8.sym # of pins=14
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/dec_3to8.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/dec_3to8.sch
.subckt dec_3to8  A1 EN A2 A0 VDD VSS Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7   NF=2
*.PININFO A2:I A1:I A0:I VDD:B VSS:B Y0:O Y1:O Y2:O Y3:O Y4:O Y5:O Y6:O Y7:O EN:I
X_inv7 A2 VDD VSS net3 inv NF=2
X_inv8 A1 VDD VSS net2 inv NF=2
X_inv9 A0 VDD VSS net1 inv NF=2
x_AndF1 net3 net2 Y0 VDD VSS net1 EN and_4in NF=1
x_AndF2 net3 net2 Y1 VDD VSS A0 EN and_4in NF=1
x_AndF3 net3 A1 Y2 VDD VSS net1 EN and_4in NF=1
x_AndF4 net3 A1 Y3 VDD VSS A0 EN and_4in NF=1
x_AndF5 A2 net2 Y4 VDD VSS net1 EN and_4in NF=1
x_AndF6 A2 net2 Y5 VDD VSS A0 EN and_4in NF=1
x_AndF7 A2 A1 Y6 VDD VSS net1 EN and_4in NF=1
x_AndF8 A2 A1 Y7 VDD VSS A0 EN and_4in NF=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/inv.sym # of pins=4
** sym_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/inv.sym
** sch_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/inv.sch
.subckt inv  X VDD VSS Y   NF=2
*.PININFO VSS:B X:I Y:O VDD:B
XM1 Y X VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y X VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/byte_dff.sym # of pins=22
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/byte_dff.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/byte_dff.sch
.subckt byte_dff  VDD VSS WE Di<3> Di<7> Do<3> Do<7> CLK SEL Di<2> Di<6> Do<2> Do<6> Di<5> Di<1>
+ Do<5> Do<1> Di<4> Do<4> Di<0> Do<0> RE   NF=2
*.PININFO Do<7>:O Di<7>:I Do<6>:O Di<6>:I Do<5>:O Di<5>:I Do<4>:O Di<4>:I Do<3>:O Di<3>:I Do<2>:O
*+ Di<2>:I Do<1>:O Di<1>:I Do<0>:O Di<0>:I WE:I SEL:I CLK:I VDD:B VSS:B RE:I
X_nand1 SEL WE net1 VDD VSS nand NF=1
X_inv1 net1 VDD VSS net2 inv NF=2
X_inv2 RE VDD VSS RE_bar inv NF=NF*3
x1 VDD net2 ck_o CLK VSS clk_gate NF=2
xDFF1 VDD VSS tinv_in7 dffout7 Di<7> ck_o DFF NF=1
X_tinv1 tinv_in7 RE_buf RE_bar VDD VSS Do<7> tinv NF=NF
xDFF2 VDD VSS tinv_in6 dffout6 Di<6> ck_o DFF NF=1
xDFF3 VDD VSS tinv_in5 dffout5 Di<5> ck_o DFF NF=1
xDFF4 VDD VSS tinv_in4 dffout4 Di<4> ck_o DFF NF=1
xDFF5 VDD VSS tinv_in3 dffout3 Di<3> ck_o DFF NF=1
xDFF6 VDD VSS tinv_in2 dffout2 Di<2> ck_o DFF NF=1
xDFF7 VDD VSS tinv_in1 dffout1 Di<1> ck_o DFF NF=1
xDFF8 VDD VSS tinv_in0 dffout0 Di<0> ck_o DFF NF=1
X_tinv2 tinv_in6 RE_buf RE_bar VDD VSS Do<6> tinv NF=NF
X_tinv3 tinv_in5 RE_buf RE_bar VDD VSS Do<5> tinv NF=NF
X_tinv4 tinv_in4 RE_buf RE_bar VDD VSS Do<4> tinv NF=NF
X_tinv5 tinv_in3 RE_buf RE_bar VDD VSS Do<3> tinv NF=NF
X_tinv6 tinv_in2 RE_buf RE_bar VDD VSS Do<2> tinv NF=NF
X_tinv7 tinv_in1 RE_buf RE_bar VDD VSS Do<1> tinv NF=NF
X_tinv8 tinv_in0 RE_buf RE_bar VDD VSS Do<0> tinv NF=NF
X_inv3 RE_bar VDD VSS RE_buf inv NF=NF*3
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/nand.sym # of pins=5
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nand.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nand.sch
.subckt nand  B A Y VDD VSS   NF=2
*.PININFO Y:O A:I VDD:B VSS:B B:I
XM2 net1 B VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y B VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 Y A VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 Y A net1 VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/and_4in.sym # of pins=7
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/and_4in.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/and_4in.sch
.subckt and_4in  A0 A1 OUT VDD VSS A2 A3   NF=1
*.PININFO VSS:B VDD:B A0:I A1:I A2:I A3:I OUT:O
X_nand1 A1 A0 net1 VDD VSS nand NF=NF
X_nand2 A3 A2 net2 VDD VSS nand NF=NF
X_nor1 OUT net1 net2 VDD VSS nor NF=NF
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/clk_gate.sym # of pins=5
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/clk_gate.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/clk_gate.sch
.subckt clk_gate  VDD EN CK_O CK_I VSS   NF=2
*.PININFO CK_I:I VDD:B VSS:B EN:I CK_O:O
X_inv1 CK_I VDD VSS net1 inv NF=NF
X_latch1 EN net1 CK_I VSS VDD net2 latch NF=NF
X_nand1 CK_I net2 net3 VDD VSS nand NF=NF
X_inv2 net3 VDD VSS CK_O inv NF=NF*3
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/DFF.sym # of pins=6
** sym_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/DFF.sym
** sch_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/DFF.sch
.subckt DFF  VDD VSS O_bar O I CLK   NF=1
*.PININFO VDD:B VSS:B I:I CLK:I O:O O_bar:O
X_latch1 I clk_bar CLK VSS VDD net1 latch NF=1
X_latch2 net1 CLK clk_bar VSS VDD net2 latch NF=1
X_inv1 CLK VDD VSS clk_bar inv NF=1
X_inv3 net2 VDD VSS O_bar inv NF=NF
X_inv4 O_bar VDD VSS O inv NF=NF
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/tinv.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv.sch
.subckt tinv  X EN ENB VDD VSS Y   NF=2
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y ENB net2 VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y EN net1 VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 X VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/nor.sym # of pins=5
** sym_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nor.sym
** sch_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nor.sch
.subckt nor  Y A B VDD VSS   NF=2
*.PININFO VDD:B VSS:B Y:O A:I B:I
XM3 net1 B VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 Y A net1 VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 Y B VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y A VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/latch.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/latch.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/latch.sch
.subckt latch  IN CLK CLKB VSS VDD OUT   NF=2
*.PININFO CLKB:I IN:I CLK:I VDD:B VSS:B OUT:O
X_tinv1 IN CLK CLKB VDD VSS net1 tinv NF=NF
X_inv1 net1 VDD VSS OUT inv NF=NF
X_tinv_small1 OUT CLKB CLK VDD VSS net1 tinv_small
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/tinv_small.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv_small.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv_small.sch
.subckt tinv_small  X EN ENB VDD VSS Y
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD pfet_03v3 L=0.28u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y ENB net2 VDD pfet_03v3 L=0.28u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y EN net1 VSS nfet_03v3 L=0.28u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 X VSS VSS nfet_03v3 L=0.28u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.end
