* NGSPICE file created from ram8_flat.ext - technology: gf180mcuC

.subckt ram8_flat A0 A1 A2 CLK Di0 Di1 Di16 Di17 Di18 Di19 Di2 Di20 Di21 Di22 Di23
+ Di24 Di25 Di26 Di27 Di28 Di29 Di3 Di30 Di31 Di4 Di5 Di6 Di7 Do0_buf Do16_buf Do17_buf
+ Do18_buf Do19_buf Do1_buf Do20_buf Do21_buf Do22_buf Do23_buf Do24_buf Do25_buf
+ Do26_buf Do27_buf Do28_buf Do29_buf Do2_buf Do30_buf Do31_buf Do3_buf Do4_buf Do5_buf
+ Do6_buf Do7_buf EN RE WE0 WE1 WE2 WE3 VSS VDD
X0 VDD a_151860_11764# a_151820_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1 a_108840_10088# a_108630_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2 word4.byte2.tinv7.O word4.byte2.tinv5.EN a_121080_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3 a_153300_306# word1.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4 VSS word6.byte4.tinv6.I a_24420_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5 VDD a_60420_9714# a_61980_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6 a_65020_6412# word5.byte3.cgate0.inv1.O a_65250_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7 Do18_buf buf_out19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8 a_124680_6578# word5.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9 word2.byte1.dff_7.O word2.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10 word7.byte1.dff_0.O word7.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11 VSS word1.byte1.cgate0.nand0.B word1.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12 VSS word2.byte4.buf_RE0.O word2.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X13 VSS word4.gt_re1.O word4.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X14 VDD word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X15 word4.byte1.cgate0.nand0.A word4.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X16 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X17 a_119430_7978# a_118810_8768# a_119320_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X18 a_15570_4842# a_14950_5632# a_15460_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X19 VDD word8.byte4.tinv2.I a_10020_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X20 word5.byte3.cgate0.nand0.A word5.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X21 a_119640_6952# a_119430_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X22 a_65020_3276# word3.byte3.cgate0.inv1.O a_65250_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X23 a_47580_5912# word4.byte3.cgate0.inv1.O a_47020_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X24 VSS a_60420_9714# a_61980_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X25 VSS word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X26 a_134580_3442# word3.byte1.cgate0.nand0.A word3.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X27 a_124680_3442# word3.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X28 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X29 VDD CLK word1.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X30 word4.byte4.dff_7.O word4.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X31 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X32 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X33 a_114880_7928# a_115210_8768# a_115110_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X34 VSS word1.byte1.cgate0.nand0.B word1.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X35 word2.byte1.cgate0.nand0.A word2.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X36 VDD word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X37 a_15570_1706# a_14950_2496# a_15460_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X38 a_119640_3816# a_119430_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X39 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X40 word3.byte3.cgate0.nand0.A word3.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X41 VDD a_153300_4840# a_154860_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X42 word4.byte2.cgate0.inv1.I word4.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X43 a_61750_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X44 a_1380_680# a_1170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X45 a_14850_2776# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X46 word8.byte3.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X47 word2.byte4.dff_7.O word2.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X48 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X49 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X50 a_140850_6462# word5.byte1.dff_7.CLK a_140740_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X51 buf_in16.inv0.O buf_in16.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X52 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X53 VDD word4.byte3.tinv3.I a_53220_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X54 a_147660_9598# word7.byte1.dff_7.CLK a_147100_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X55 VDD a_100380_6462# a_101040_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X56 VDD a_153300_1704# a_154860_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X57 word2.byte2.cgate0.inv1.I word2.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X58 a_47970_9598# word7.byte3.cgate0.inv1.O a_47860_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X59 a_61750_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X60 VDD buf_in9.inv0.O buf_in9.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X61 VSS word8.byte2.tinv4.I a_117480_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X62 a_140130_9598# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X63 VDD word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X64 a_24420_6578# word5.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X65 VDD a_42420_306# a_43980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X66 a_140850_3326# word3.byte1.dff_7.CLK a_140740_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X67 word7.byte3.dff_5.O word7.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X68 word7.byte4.tinv7.O buf_out30.inv0.I a_10020_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X69 a_111610_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X70 VSS a_166260_8628# a_166220_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X71 VDD word2.byte3.tinv3.I a_53220_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X72 VSS buf_in28.inv0.O buf_in28.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X73 VDD a_100380_3326# a_101040_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X74 a_155140_4842# a_153300_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X75 VSS a_110280_1704# a_111840_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X76 VDD a_55380_5492# a_55340_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X77 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X78 VSS word2.byte1.tinv0.I a_142500_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X79 a_142500_11112# word8.byte1.tinv0.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X80 a_19380_680# a_19170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X81 VDD word5.byte4.dff_0.O_bar a_2820_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X82 VSS a_1380_680# word1.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X83 a_155140_1706# a_153300_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X84 a_48140_9598# a_47350_9548# a_47970_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X85 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X86 a_122410_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X87 VSS word2.byte2.inv_and.O a_92280_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X88 VDD a_55380_2356# a_55340_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X89 a_4770_7978# word6.byte4.cgate0.inv1.O a_4660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X90 a_123030_4842# word4.byte2.dff_7.CLK a_122920_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X91 VSS word8.byte4.dff_0.O_bar a_2820_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X92 VDD EN dec8.and4_1.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X93 word6.byte2.dff_2.O word6.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X94 VDD word3.byte4.dff_0.O_bar a_2820_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X95 a_131700_9714# word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X96 a_156900_11112# buf_out4.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X97 VSS a_162660_680# a_162620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X98 VSS word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X99 VSS word1.byte4.tinv5.I a_20820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X100 word5.byte1.nand.B word5.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X101 VSS word8.gt_re0.OUT word8.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X102 a_11860_10498# a_10020_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X103 word7.byte2.cgate0.nand0.A word7.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X104 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X105 a_54780_2776# word2.byte3.cgate0.inv1.O a_54220_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X106 word5.byte3.tinv7.O buf_out23.inv0.I a_46020_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X107 VSS a_108840_680# a_108800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X108 word3.byte1.nand.B word3.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X109 VSS buf_out13.inv0.I buf_out13.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X110 a_25980_9048# word6.byte4.cgate0.inv1.O a_25420_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X111 a_54450_11114# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X112 a_108240_12184# word8.byte2.dff_7.CLK a_107680_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X113 word3.byte3.tinv7.O buf_out23.inv0.I a_46020_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X114 a_65860_5912# a_64020_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X115 a_13620_4840# word4.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X116 a_119600_11114# word8.byte2.dff_7.CLK a_119430_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X117 a_159020_10498# word7.byte1.dff_7.CLK a_158850_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X118 VDD word8.buf_ck1.I word8.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X119 a_50850_6462# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X120 VSS buf_in6.inv0.O buf_in6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X121 a_40770_190# word1.byte3.cgate0.inv1.O a_40660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X122 a_7980_1090# a_7750_140# a_7420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X123 a_161730_7362# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X124 a_13620_1704# word2.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X125 VDD buf_out24.inv0.I buf_out24.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X126 buf_we4.inv1.O buf_we4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X127 a_22660_7978# a_20820_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X128 a_50850_3326# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X129 VSS word6.buf_sel0.O word6.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X130 a_66180_5492# a_65970_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X131 a_108840_2356# a_108630_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X132 a_161730_4226# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X133 VSS buf_out31.inv0.I buf_out31.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X134 a_165660_10498# a_165430_9548# a_165100_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X135 a_162060_1090# a_161830_140# a_161500_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X136 a_62370_190# a_61750_140# a_62260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X137 a_118810_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X138 a_155250_4842# word4.byte1.dff_7.CLK a_155140_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X139 a_101600_5912# a_100810_5632# a_101430_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X140 buf_in21.inv1.O buf_in21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X141 a_4940_11114# word8.byte4.cgate0.inv1.O a_4770_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X142 a_53220_11112# word8.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X143 a_100710_4842# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X144 word1.byte1.dff_3.O word1.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X145 word2.byte3.tinv7.O word2.byte3.tinv6.EN a_64020_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X146 VSS a_19380_5492# word4.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X147 a_22980_8628# a_22770_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X148 buf_sel3.inv1.O buf_sel3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X149 a_107680_11064# word8.byte2.dff_7.CLK a_107910_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X150 a_147100_9548# word7.byte1.dff_7.CLK a_147330_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X151 a_166260_10088# a_166050_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X152 word1.byte1.tinv7.O buf_out2.inv0.I a_164100_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X153 VDD a_53220_11112# a_54780_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X154 VDD word1.byte2.tinv2.I a_110280_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X155 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X156 VSS a_66180_2356# word2.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X157 a_65350_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X158 a_100710_1706# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X159 a_167700_4840# buf_out1.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X160 a_119600_9048# a_118810_8768# a_119430_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X161 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X162 VSS word7.byte3.dff_0.O_bar a_42420_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X163 a_35760_3442# word3.byte1.cgate0.nand0.B word3.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X164 VSS word5.byte1.buf_RE1.I word5.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X165 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X166 a_67620_11112# word8.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X167 a_62540_7978# word6.byte3.cgate0.inv1.O a_62370_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X168 a_167700_1704# buf_out1.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X169 VDD word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X170 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X171 word5.byte1.nand.B word5.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X172 a_75720_4840# word4.byte3.cgate0.latch0.I0.ENB word4.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X173 a_62260_7362# a_60420_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X174 VSS a_100380_11114# a_101040_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X175 word1.buf_sel0.O buf_sel1.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X176 a_148260_680# a_148050_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X177 a_139900_6412# a_140230_6412# a_140130_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X178 VDD a_147100_9548# a_146100_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X179 buf_in12.inv0.O buf_in12.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X180 a_56820_7976# buf_out20.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X181 VDD a_112440_11764# a_112400_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X182 VDD a_151860_10088# a_151820_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X183 a_47350_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X184 a_115210_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X185 a_75720_1704# word2.byte3.cgate0.latch0.I0.ENB word2.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X186 a_450_4842# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X187 buf_in3.inv0.O Di2 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X188 a_65970_190# word1.byte3.cgate0.inv1.O a_65860_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X189 a_62260_4226# a_60420_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X190 VSS buf_out26.inv0.O Do25_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X191 a_139900_3276# a_140230_3276# a_140130_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X192 VDD a_162660_6952# word5.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X193 a_62580_6952# a_62370_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X194 VDD buf_out8.inv0.O Do7_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X195 VDD buf_out29.inv0.I buf_out29.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X196 a_450_1706# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X197 a_146100_4840# word4.byte1.tinv1.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X198 a_8370_7978# a_7750_8768# a_8260_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X199 a_7420_140# a_7750_140# a_7650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X200 VDD a_162660_3816# word3.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X201 word4.byte1.dff_1.O word4.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X202 Do17_buf buf_out18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X203 VSS word6.byte3.tinv2.I a_49620_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X204 a_62580_3816# a_62370_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X205 word2.byte1.cgate0.inv1.I word2.byte1.cgate0.nand0.A a_134580_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X206 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X207 buf_in32.inv0.O Di31 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X208 a_122080_4792# a_122410_5632# a_122310_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X209 VDD word5.byte1.tinv2.I a_149700_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X210 VSS word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X211 VDD a_101640_5492# word4.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X212 word8.byte2.dff_7.O word8.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X213 VSS word3.byte1.tinv5.I a_160500_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X214 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X215 a_106680_6578# buf_out15.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X216 a_162450_1706# word2.byte1.dff_7.CLK a_162340_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X217 VSS a_26580_6952# a_26540_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X218 VDD word3.byte1.tinv2.I a_149700_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X219 VDD a_101640_2356# word2.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X220 a_65250_5912# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X221 VDD buf_sel1.inv0.I buf_sel1.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X222 a_11020_140# word1.byte4.cgate0.inv1.O a_11250_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X223 VSS word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X224 word3.byte2.tinv7.O word3.byte2.tinv4.EN a_117480_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X225 a_106680_3442# buf_out15.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X226 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X227 VSS a_108840_11764# word8.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X228 a_40050_2776# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X229 VSS word3.byte1.nand.OUT word3.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X230 VDD word5.byte3.buf_RE0.O word5.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X231 VSS a_26580_3816# a_26540_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X232 a_166050_6462# word5.byte1.dff_7.CLK a_165940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X233 a_106680_9714# word7.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X234 VSS buf_in15.inv0.O buf_in15.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X235 VDD a_147100_7928# a_146100_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X236 VDD a_124680_6578# a_126240_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X237 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X238 word4.byte2.inv_and.O word4.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X239 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X240 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X241 a_165330_9598# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X242 a_49620_6578# word5.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X243 VDD word3.byte3.buf_RE0.O word3.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X244 VDD buf_out9.inv0.I buf_out9.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X245 a_166050_3326# word3.byte1.dff_7.CLK a_165940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X246 word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.latch0.I0.ENB a_36120_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X247 VDD word6.byte1.nand.B word6.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X248 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.latch0.I0.ENB a_131700_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X249 word2.byte2.inv_and.O word2.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X250 VDD a_124680_3442# a_126240_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X251 a_108520_5912# a_106680_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X252 word6.byte4.tinv7.O buf_out28.inv0.I a_17220_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X253 VDD a_119640_11764# word8.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X254 VSS word2.byte1.tinv7.I a_167700_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X255 word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.latch0.I0.ENB a_36120_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X256 VDD buf_in11.inv0.I buf_in11.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X257 VDD buf_in25.inv0.O buf_in25.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X258 VDD a_116040_680# word1.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X259 word5.byte1.dff_0.O word5.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X260 a_22940_12184# a_22150_11904# a_22770_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X261 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.latch0.I0.O a_131700_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X262 VDD a_61420_6412# a_60420_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X263 a_124680_1704# word2.byte2.tinv6.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X264 VSS Di1 buf_in2.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X265 a_48140_12184# a_47350_11904# a_47970_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X266 a_117480_11112# buf_out12.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X267 a_147330_1090# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X268 a_69420_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X269 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X270 a_75360_2660# word2.byte1.cgate0.nand0.B word2.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X271 VSS a_108840_10088# a_108800_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X272 word6.gt_re0.OUT buf_sel6.inv1.O a_82020_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X273 a_50620_6412# word5.byte3.cgate0.inv1.O a_50850_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X274 VSS a_15780_680# a_15740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X275 word3.byte1.dff_0.O word3.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X276 VDD buf_in31.inv0.O buf_in31.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X277 buf_in19.inv1.O buf_in19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X278 word2.byte1.dff_3.O word2.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X279 VDD a_61420_3276# a_60420_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X280 a_156900_9714# word7.byte1.tinv4.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X281 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X282 VSS word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X283 VSS word4.byte3.tinv4.I a_56820_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X284 VDD word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X285 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X286 a_105030_7978# a_104410_8768# a_104920_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X287 a_50620_3276# word3.byte3.cgate0.inv1.O a_50850_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X288 buf_sel2.inv1.O buf_sel2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X289 a_54450_10498# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X290 a_6420_7976# word6.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X291 a_100480_7928# a_100810_8768# a_100710_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X292 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X293 a_2820_11112# buf_out32.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X294 a_119600_10498# word7.byte2.dff_7.CLK a_119430_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X295 word4.byte1.tinv7.O buf_out3.inv0.I a_160500_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X296 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X297 a_11020_11064# a_11350_11904# a_11250_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X298 word7.byte3.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X299 word3.gt_re1.O word3.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X300 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X301 VDD word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X302 a_54550_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X303 a_150930_11114# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X304 a_151030_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X305 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X306 a_144620_6462# a_143830_6412# a_144450_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X307 a_22770_11114# a_22150_11904# a_22660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X308 a_43650_9048# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X309 VDD a_57820_4792# a_56820_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X310 VDD buf_out15.inv0.O buf_out15.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X311 word7.byte2.dff_3.O word7.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X312 VSS a_166260_10088# word7.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X313 word2.byte1.tinv7.O buf_out3.inv0.I a_160500_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X314 VSS word3.byte4.tinv7.I a_28020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X315 buf_in32.inv1.O buf_in32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X316 VDD word8.gt_re1.O word8.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X317 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X318 VDD word7.byte2.tinv2.I a_110280_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X319 VSS a_151860_8628# a_151820_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X320 VSS buf_out6.inv0.O Do5_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X321 a_144620_3326# a_143830_3276# a_144450_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X322 a_140740_4842# a_139800_4842# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X323 VDD a_57820_1656# a_56820_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X324 VDD a_40980_5492# a_40940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X325 VDD a_139900_11064# a_139800_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X326 word6.byte3.tinv7.O buf_out22.inv0.I a_49620_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X327 a_159060_5492# a_158850_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X328 VDD buf_re.inv0.O buf_re.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X329 a_115720_2776# a_113880_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X330 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X331 a_40980_11764# a_40770_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X332 a_4940_10498# word7.byte4.cgate0.inv1.O a_4770_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X333 a_47860_7978# a_46020_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X334 a_58150_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X335 a_140740_1706# a_139800_1706# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X336 a_220_7928# a_550_8768# a_450_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X337 VSS word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X338 VDD a_40980_2356# a_40940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X339 buf_in20.inv1.O buf_in20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X340 a_107680_9548# word7.byte2.dff_7.CLK a_107910_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X341 a_159060_2356# a_158850_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X342 VDD a_148260_680# word1.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X343 VDD a_53220_9714# a_54780_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X344 a_58150_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X345 a_126800_5912# a_126010_5632# a_126630_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X346 a_7420_1656# a_7750_2496# a_7650_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X347 a_125910_4842# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X348 VSS a_44580_5492# word4.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X349 a_42420_7976# word6.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X350 VSS a_61420_7928# a_60420_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X351 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X352 a_48180_8628# a_47970_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X353 dec8.and4_5.nand0.OUT A0 a_73020_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X354 a_142500_6578# word5.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X355 VDD word8.byte4.tinv7.I a_28020_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X356 a_125910_1706# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X357 VSS word4.buf_sel0.O word4.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X358 a_15740_1090# word1.byte4.cgate0.inv1.O a_15570_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X359 a_164100_6578# word5.byte1.tinv6.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X360 buf_sel8.inv1.O buf_sel8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X361 a_92280_7364# word5.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X362 VDD word5.byte2.buf_RE1.I word5.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X363 VSS word7.byte3.tinv7.I a_67620_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X364 VSS a_24420_6578# a_25980_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X365 a_142500_3442# word3.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X366 VDD a_112440_10088# a_112400_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X367 word1.byte2.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B a_93540_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X368 VDD a_123240_680# a_123200_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X369 VSS a_148260_680# word1.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X370 VSS word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X371 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X372 VDD word3.byte2.buf_RE1.I word3.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X373 a_92280_4228# word3.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X374 a_21820_4792# word4.byte4.cgate0.inv1.O a_22050_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X375 VSS a_24420_3442# a_25980_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X376 a_165100_6412# a_165430_6412# a_165330_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X377 VSS word5.byte4.buf_RE0.O word5.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X378 VSS a_146100_1704# a_147660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X379 VDD word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X380 a_122920_190# a_121080_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X381 a_21820_1656# word2.byte4.cgate0.inv1.O a_22050_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X382 buf_out11.inv1.O buf_out11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X383 word7.byte4.tinv7.O buf_out25.inv0.I a_28020_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X384 VSS a_65020_9548# a_64020_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X385 a_165100_3276# a_165430_3276# a_165330_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X386 VDD buf_in7.inv0.O buf_in7.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X387 VDD word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X388 a_119640_5492# a_119430_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X389 a_158460_190# word1.byte1.dff_7.CLK a_157900_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X390 a_54220_9548# a_54550_9548# a_54450_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X391 a_160500_1704# word2.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X392 a_161830_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X393 buf_in31.inv0.O Di30 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X394 VDD a_104080_6412# a_103080_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X395 a_123200_7362# word5.byte2.dff_7.CLK a_123030_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X396 VSS a_48180_2356# a_48140_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X397 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X398 a_33420_12068# word8.byte4.cgate0.nand0.A word8.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X399 VDD a_126840_5492# word4.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X400 a_140850_4842# word4.byte1.dff_7.CLK a_140740_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X401 Do21_buf buf_out22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X402 VSS a_55380_11764# word8.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X403 a_132960_7364# word5.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X404 a_161830_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X405 VSS a_19380_8628# a_19340_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X406 VDD a_47020_140# a_46020_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X407 VSS CLK word4.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X408 a_123200_4226# word3.byte2.dff_7.CLK a_123030_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X409 VDD a_104080_3276# a_103080_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X410 buf_sel2.inv1.O buf_sel2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X411 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X412 a_158130_4842# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X413 VSS a_51780_2356# word2.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X414 VSS word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X415 VDD a_126840_2356# word2.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X416 a_50950_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X417 word7.byte1.tinv7.O word7.byte1.tinv2.EN a_149700_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X418 a_132960_4228# word3.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X419 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X420 VDD A1 dec8.and4_6.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X421 a_104080_7928# word6.byte2.dff_7.CLK a_104310_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X422 a_158850_7978# word6.byte1.dff_7.CLK a_158740_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X423 VSS a_22980_8628# word6.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X424 a_158130_1706# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X425 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X426 VDD word6.byte1.tinv3.I a_153300_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X427 a_28020_9714# word7.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X428 VDD a_21820_11064# a_20820_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X429 a_144340_11114# a_142500_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X430 a_56820_306# buf_out20.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X431 VDD a_47020_11064# a_46020_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X432 VSS word8.byte2.inv_and.O a_92280_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X433 VDD a_119640_10088# word7.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X434 a_47250_7978# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X435 a_110280_7976# buf_out14.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X436 VDD word5.byte4.tinv2.I a_10020_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X437 VDD a_4980_680# word1.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X438 word4.byte3.cgate0.inv1.I word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X439 VDD buf_in12.inv0.O buf_in12.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X440 VSS word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X441 VDD word8.byte1.cgate0.nand0.B word8.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X442 a_100810_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X443 VDD a_155460_8628# a_155420_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X444 a_141020_190# a_140230_140# a_140850_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X445 a_144060_6462# word5.byte1.dff_7.CLK a_143500_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X446 a_44370_6462# word5.byte3.cgate0.inv1.O a_44260_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X447 VDD word3.byte4.tinv2.I a_10020_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X448 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X449 VSS a_149700_7976# a_151260_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X450 word5.byte3.dff_4.O word5.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X451 word2.byte3.cgate0.inv1.I word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X452 buf_in10.inv1.O buf_in10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X453 VDD buf_in6.inv0.O buf_in6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X454 a_144060_3326# word3.byte1.dff_7.CLK a_143500_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X455 VDD a_39720_4842# a_40380_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X456 word6.byte1.tinv7.O word6.byte1.tinv4.EN a_156900_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X457 a_44370_3326# word3.byte3.cgate0.inv1.O a_44260_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X458 word5.byte1.dff_7.O word5.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X459 VSS word6.byte2.tinv0.I a_103080_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X460 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X461 a_111840_11114# a_111610_11904# a_111280_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X462 a_144620_12184# a_143830_11904# a_144450_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X463 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X464 VDD word7.byte1.tinv7.I a_167700_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X465 buf_we2.inv0.O WE1 VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X466 buf_in1.inv1.O buf_in1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X467 word3.byte3.dff_4.O word3.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X468 word6.byte4.dff_1.O word6.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X469 a_46020_11112# word8.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X470 VDD a_39720_1706# a_40380_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X471 word3.byte1.dff_7.O word3.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X472 VDD buf_in30.inv0.O buf_in30.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X473 Do26_buf buf_out27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X474 VSS word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X475 a_14850_7362# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X476 word4.byte2.dff_1.O word4.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X477 VSS A0 dec8.and4_6.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X478 VSS a_104080_7928# a_103080_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X479 word6.byte1.dff_5.O word6.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X480 a_151260_12184# word8.byte1.dff_7.CLK a_150700_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X481 VSS a_143500_140# a_142500_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X482 a_50850_5912# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X483 buf_sel3.inv1.O buf_sel3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X484 VSS word8.byte1.nand.B a_78780_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X485 a_111510_11114# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X486 a_150930_10498# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X487 a_166220_2776# a_165430_2496# a_166050_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X488 a_22770_9598# a_22150_9548# a_22660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X489 VSS a_47020_1656# a_46020_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X490 word2.byte2.dff_1.O word2.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X491 word3.byte2.tinv7.O word3.byte2.tinv0.EN a_103080_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X492 a_95160_3442# word3.byte2.cgate0.nand0.A word3.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X493 a_14850_4226# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X494 a_15180_1090# a_14950_140# a_14620_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X495 a_60420_9714# word7.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X496 a_95160_6578# word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X497 a_103080_6578# word5.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X498 VDD a_110280_6578# a_111840_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X499 a_26540_4842# word4.byte4.cgate0.inv1.O a_26370_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X500 VDD a_139900_9548# a_139800_9598# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X501 VDD word1.byte1.nand.B word1.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X502 a_4660_2776# a_2820_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X503 VSS a_117480_11112# a_119040_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X504 a_150930_9598# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X505 a_40980_10088# a_40770_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X506 word1.byte4.tinv7.O buf_out28.inv0.I a_17220_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X507 a_19380_10088# a_19170_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X508 a_126240_9048# word6.byte2.dff_7.CLK a_125680_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X509 VDD a_53220_306# a_54780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X510 VSS a_160500_306# a_162060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X511 a_26540_1706# word2.byte4.cgate0.inv1.O a_26370_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X512 VDD a_110280_3442# a_111840_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X513 VSS buf_out28.inv0.O Do27_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X514 VDD word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X515 a_165940_4842# a_164100_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X516 VDD word6.byte3.cgate0.nand0.A a_75360_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X517 a_110280_11112# word8.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X518 a_162660_11764# a_162450_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X519 a_4980_2356# a_4770_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X520 a_58940_9598# a_58150_9548# a_58770_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X521 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X522 a_165940_1706# a_164100_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X523 Do19_buf buf_out20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X524 a_115110_190# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X525 word4.byte1.tinv7.O word4.byte1.tinv6.EN a_164100_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X526 VSS word4.byte2.tinv2.I a_110280_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X527 a_67620_8932# word6.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X528 a_54780_7362# a_54550_6412# a_54220_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X529 a_4150_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X530 a_139900_4792# a_140230_5632# a_140130_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X531 a_167700_7364# word5.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X532 a_124680_11112# word8.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X533 a_6420_306# word1.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X534 a_160500_306# word1.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X535 a_24420_7976# word6.byte4.tinv6.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X536 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X537 VSS word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X538 a_108800_7978# word6.byte2.dff_7.CLK a_108630_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X539 word5.byte2.tinv7.O buf_out10.inv0.I a_124680_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X540 buf_we3.inv1.O buf_we3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X541 a_162660_6952# a_162450_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X542 VDD a_26580_8628# word6.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X543 a_167700_4228# word3.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X544 a_54780_4226# a_54550_3276# a_54220_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X545 VSS a_111280_4792# a_110280_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X546 a_51460_9598# a_49620_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X547 word4.byte1.cgate0.inv1.I word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X548 word8.byte1.tinv7.O buf_out6.inv0.I a_149700_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X549 a_157900_7928# a_158230_8768# a_158130_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X550 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X551 a_106680_306# word1.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X552 word3.byte2.tinv7.O buf_out10.inv0.I a_124680_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X553 a_162660_3816# a_162450_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X554 a_47020_4792# word4.byte3.cgate0.inv1.O a_47250_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X555 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X556 VDD word4.gt_re1.O word4.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X557 VDD buf_sel5.inv0.O buf_sel5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X558 word2.byte1.cgate0.inv1.I word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X559 VSS word3.byte4.tinv3.I a_13620_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X560 VDD buf_in15.inv0.O buf_in15.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X561 VSS a_151860_10088# word7.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X562 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X563 word1.byte3.tinv7.O buf_out22.inv0.I a_49620_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X564 word8.byte1.nand.B word8.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X565 a_51780_10088# a_51570_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X566 a_47020_1656# word2.byte3.cgate0.inv1.O a_47250_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X567 a_108840_6952# a_108630_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X568 VDD word2.gt_re1.O word2.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X569 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X570 VSS buf_in6.inv0.O buf_in6.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X571 a_53220_4840# buf_out21.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X572 a_154630_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X573 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X574 word5.byte4.tinv7.O word5.byte4.tinv6.EN a_24420_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X575 VSS a_26580_5492# a_26540_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X576 a_43750_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X577 a_108840_3816# a_108630_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X578 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X579 a_53220_1704# buf_out21.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X580 VSS buf_in30.inv0.O buf_in30.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X581 a_10020_9714# word7.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X582 Do26_buf buf_out27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X583 VDD a_66180_6952# word5.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X584 VSS a_117480_306# a_119040_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X585 a_18450_9598# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X586 a_142500_1704# word2.byte1.tinv0.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X587 a_43750_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X588 a_166050_4842# word4.byte1.dff_7.CLK a_165940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X589 buf_in21.inv1.O buf_in21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X590 Do1_buf buf_out2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X591 a_6420_11112# word8.byte4.tinv1.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X592 a_101640_8628# a_101430_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X593 a_2820_6578# buf_out32.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X594 a_92280_2660# word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X595 VSS buf_out19.inv0.O Do18_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X596 VDD a_66180_3816# word3.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X597 a_47580_12184# word8.byte3.cgate0.inv1.O a_47020_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X598 VSS word7.byte2.tinv5.I a_121080_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X599 a_2820_3442# buf_out32.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X600 buf_sel8.inv0.I dec8.and4_7.nand1.OUT a_77700_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X601 a_51740_11114# word8.byte3.cgate0.inv1.O a_51570_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X602 a_144340_10498# a_142500_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X603 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X604 VSS a_10020_6578# a_11580_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X605 VSS a_113880_9714# a_115440_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X606 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X607 VSS a_161500_6412# a_160500_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X608 VDD word7.buf_ck1.I word7.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X609 a_7650_6462# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X610 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X611 VDD a_143500_11064# a_142500_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X612 VSS a_10020_3442# a_11580_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X613 VDD word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X614 a_126010_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X615 VSS a_161500_3276# a_160500_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X616 word6.byte3.dff_2.O word6.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X617 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X618 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X619 a_7650_3326# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X620 a_105200_12184# a_104410_11904# a_105030_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X621 buf_in9.inv1.O buf_in9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X622 a_50950_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X623 a_111840_10498# a_111610_9548# a_111280_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X624 VDD word7.byte2.tinv7.I a_128280_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X625 VSS a_50620_9548# a_49620_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X626 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X627 VSS word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X628 VSS word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X629 VDD buf_in28.inv0.O buf_in28.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X630 a_58980_11764# a_58770_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X631 VDD a_64020_4840# a_65580_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X632 word4.byte4.tinv7.O buf_out29.inv0.I a_13620_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X633 a_39820_11064# word8.byte3.cgate0.inv1.O a_40050_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X634 VSS word6.byte2.tinv7.I a_128280_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X635 word2.byte1.cgate0.nand0.A word2.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X636 a_92280_11112# word8.byte2.cgate0.latch0.I0.ENB word8.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X637 VDD word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X638 a_153300_9714# buf_out5.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X639 VSS a_4980_10088# a_4940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X640 Do25_buf buf_out26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X641 a_58380_9598# word7.byte3.cgate0.inv1.O a_57820_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X642 a_162450_6462# a_161830_6412# a_162340_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X643 VDD a_64020_1704# a_65580_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X644 word2.byte4.tinv7.O buf_out29.inv0.I a_13620_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X645 buf_in26.inv1.O buf_in26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X646 VSS word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X647 a_167700_12068# word8.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X648 a_123240_8628# a_123030_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X649 buf_in20.inv1.O buf_in20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X650 a_111510_10498# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X651 word2.byte2.cgate0.inv1.I word2.byte2.cgate0.nand0.A a_95160_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X652 VSS a_105240_6952# a_105200_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X653 a_40050_7362# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X654 a_162450_3326# a_161830_3276# a_162340_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X655 a_144620_5912# a_143830_5632# a_144450_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X656 dec8.and4_1.nand0.OUT A0 a_65820_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X657 a_143730_4842# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X658 VSS word2.byte3.tinv3.I a_53220_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X659 VSS a_39720_11114# a_40380_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X660 a_118710_2776# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X661 a_101430_4842# a_100810_5632# a_101320_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X662 VDD word1.byte1.tinv3.I a_153300_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X663 VSS a_105240_3816# a_105200_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X664 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X665 word3.byte2.tinv7.O word3.byte2.tinv7.EN a_128280_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X666 a_40050_4226# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X667 VSS word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X668 a_143730_1706# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X669 word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.latch0.I0.O a_93540_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X670 VSS buf_sel5.inv0.O buf_sel5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X671 word8.byte3.tinv7.O buf_out23.inv0.I a_46020_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X672 a_110280_306# buf_out14.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X673 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X674 a_101430_1706# a_100810_2496# a_101320_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X675 VSS word3.byte2.nand.OUT word3.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X676 a_78780_3442# buf_we2.inv1.O word3.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X677 VSS word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X678 VDD word6.byte1.buf_RE1.I word6.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X679 VDD a_157900_7928# a_156900_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X680 VDD word5.byte1.cgate0.nand0.B word5.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X681 VSS a_13620_306# a_15180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X682 a_128280_6578# word5.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X683 buf_sel1.inv0.O buf_sel1.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X684 VDD a_141060_680# a_141020_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X685 a_36120_3442# word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X686 a_42420_9714# word7.byte3.tinv0.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X687 a_162660_10088# a_162450_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X688 word5.byte3.inv_and.O word5.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X689 word5.byte2.nand.OUT buf_we3.inv1.O a_90120_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X690 VDD CLK word8.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X691 VDD word3.byte1.cgate0.nand0.B word3.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X692 VDD a_220_7928# a_120_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X693 a_158230_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X694 word5.byte3.dff_0.O word5.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X695 word1.byte2.cgate0.inv1.I word1.byte2.cgate0.nand0.A a_95160_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X696 word5.byte1.dff_3.O word5.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X697 a_55060_190# a_53220_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X698 VSS buf_we4.inv0.O buf_we4.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X699 word3.byte3.dff_0.O word3.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X700 a_44260_4842# a_42420_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X701 VSS a_24420_4840# a_25980_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X702 a_18220_6412# a_18550_6412# a_18450_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X703 word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.latch0.I0.O a_92280_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X704 a_13620_306# word1.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X705 word3.byte1.dff_3.O word3.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X706 VDD buf_out31.inv0.O Do30_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X707 buf_in4.inv1.O buf_in4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X708 a_115830_190# a_115210_140# a_115720_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X709 a_11350_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X710 word6.byte4.inv_and.O word6.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X711 a_44260_1706# a_42420_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X712 VSS a_25420_11064# a_24420_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X713 a_18220_3276# a_18550_3276# a_18450_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X714 a_165100_4792# a_165430_5632# a_165330_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X715 VDD a_144660_5492# word4.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X716 a_15180_11114# a_14950_11904# a_14620_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X717 a_44580_5492# a_44370_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X718 VSS word8.byte1.cgate0.nand0.B word8.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X719 VSS word5.byte4.tinv1.I a_6420_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X720 a_151820_2776# a_151030_2496# a_151650_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X721 a_14950_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X722 a_13620_1704# word2.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X723 VDD a_144660_2356# word2.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X724 a_160500_3442# word3.byte1.tinv5.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X725 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X726 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X727 a_44580_2356# a_44370_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X728 a_122310_9048# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X729 a_33420_9714# word7.byte4.cgate0.nand0.A word7.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X730 a_117480_4840# word4.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X731 VSS word5.buf_ck1.I word5.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X732 a_14950_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X733 a_161830_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X734 VDD buf_sel6.inv0.O buf_sel6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X735 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X736 VDD buf_in14.inv0.O buf_in14.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X737 a_15460_12184# a_13620_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X738 a_47250_190# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X739 VDD word4.byte1.nand.B word4.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X740 a_115720_7362# a_113880_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X741 a_111840_9048# word6.byte2.dff_7.CLK a_111280_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X742 VDD word1.byte3.cgate0.nand0.A a_75360_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X743 a_49620_11112# buf_out22.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X744 a_153300_306# word1.byte1.tinv3.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X745 a_117480_1704# word2.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X746 VSS buf_in12.inv0.I buf_in12.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X747 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X748 a_49620_6578# word5.byte3.tinv2.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X749 a_58660_1090# a_56820_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X750 VDD word2.byte1.nand.B word2.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X751 a_115720_4226# a_113880_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X752 a_112400_9598# a_111610_9548# a_112230_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X753 a_7420_6412# word5.byte4.cgate0.inv1.O a_7650_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X754 word8.gt_re3.I word8.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X755 Do7_buf buf_out8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X756 VDD a_106680_4840# a_108240_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X757 buf_in20.inv1.O buf_in20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X758 VDD a_159060_680# word1.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X759 a_167700_2660# word2.byte1.tinv7.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X760 a_58980_680# a_58770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X761 a_121080_7976# word6.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X762 a_126840_8628# a_126630_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X763 a_7420_3276# word3.byte4.cgate0.inv1.O a_7650_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X764 VSS a_2820_9714# a_4380_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X765 VDD Di22 buf_in23.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X766 a_51740_10498# word7.byte3.cgate0.inv1.O a_51570_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X767 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B a_132960_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X768 VDD a_106680_1704# a_108240_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X769 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X770 a_10020_7976# word6.byte4.tinv2.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X771 VDD a_12180_680# word1.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X772 a_75720_2660# word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X773 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X774 VSS a_22980_680# a_22940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X775 a_144060_5912# word4.byte1.dff_7.CLK a_143500_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X776 a_148050_7978# a_147430_8768# a_147940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X777 word5.byte2.tinv7.O buf_out14.inv0.I a_110280_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X778 a_44370_4842# word4.byte3.cgate0.inv1.O a_44260_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X779 dec8.and4_0.nand0.OUT dec8.and4_6.nand0.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X780 a_56820_4840# word4.byte3.tinv4.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X781 word8.byte4.dff_4.O word8.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X782 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X783 VDD word7.gt_re1.O word7.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X784 word4.byte3.dff_4.O word4.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X785 VDD a_146100_6578# a_147660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X786 a_36120_11112# word8.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X787 a_143500_7928# a_143830_8768# a_143730_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X788 VSS a_123240_8628# word6.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X789 word3.byte2.tinv7.O buf_out14.inv0.I a_110280_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X790 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X791 a_155250_11114# a_154630_11904# a_155140_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X792 word6.byte4.tinv7.O buf_out31.inv0.I a_6420_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X793 VDD a_146100_3442# a_147660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X794 VDD buf_re.inv1.O word4.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X795 VDD word4.byte3.buf_RE0.O word4.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X796 a_58980_10088# a_58770_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X797 a_39820_9548# word7.byte3.cgate0.inv1.O a_40050_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X798 word6.byte4.dff_3.O word6.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X799 word7.byte1.dff_4.O word7.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X800 a_61750_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X801 a_19340_2776# a_18550_2496# a_19170_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X802 VDD word6.byte3.buf_RE0.O word6.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X803 VDD a_48180_6952# a_48140_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X804 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X805 VDD a_139800_7978# a_140460_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X806 VDD buf_re.inv1.O word2.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X807 VDD word2.byte3.buf_RE0.O word2.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X808 buf_in13.inv1.O buf_in13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X809 a_155460_11764# a_155250_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X810 word5.byte4.tinv7.O word5.byte4.tinv2.EN a_10020_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X811 a_128280_12068# word8.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X812 word8.byte2.cgate0.inv1.I word8.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X813 buf_in4.inv1.O buf_in4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X814 a_158740_2776# a_156900_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X815 VDD a_48180_3816# a_48140_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X816 buf_in25.inv1.O buf_in25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X817 VDD a_121080_11112# a_122640_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X818 VSS a_155460_11764# a_155420_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X819 VSS a_58980_2356# a_58940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X820 VDD a_114880_6412# a_113880_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X821 VDD a_15780_11764# word8.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X822 VDD a_51780_6952# word5.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X823 buf_in7.inv1.O buf_in7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X824 VDD a_57820_140# a_56820_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X825 a_140460_190# word1.byte1.dff_7.CLK a_139900_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X826 a_73020_8932# word6.byte3.cgate0.nand0.A word6.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X827 word4.byte4.dff_0.O word4.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X828 VDD a_114880_3276# a_113880_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X829 VSS buf_in19.inv0.O buf_in19.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X830 a_114880_140# word1.byte2.dff_7.CLK a_115110_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X831 VDD a_51780_3816# word3.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X832 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X833 word2.byte2.inv_and.O word2.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X834 VSS a_147100_4792# a_146100_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X835 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X836 VSS word1.byte3.tinv6.I a_64020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X837 VSS a_160500_11112# a_162060_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X838 a_126630_4842# a_126010_5632# a_126520_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X839 VSS word8.byte3.tinv7.I a_67620_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X840 VSS word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X841 word2.byte4.dff_0.O word2.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X842 VDD word5.byte1.cgate0.nand0.B word5.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X843 word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.latch0.I0.O a_36120_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X844 a_123030_11114# word8.byte2.dff_7.CLK a_122920_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X845 VSS word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X846 a_106680_9714# word7.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X847 word6.byte3.tinv7.O word6.byte3.tinv0.EN a_42420_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X848 word1.byte2.dff_4.O word1.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X849 a_90120_5796# word4.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X850 word8.byte1.tinv7.O buf_out1.inv0.I a_167700_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X851 word5.byte1.tinv7.O buf_out8.inv0.I a_142500_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X852 VDD word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X853 a_151260_2776# word2.byte1.dff_7.CLK a_150700_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X854 VSS buf_sel2.inv0.O buf_sel2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X855 a_119320_9598# a_117480_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X856 a_15460_6462# a_13620_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X857 a_51570_1706# word2.byte3.cgate0.inv1.O a_51460_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X858 a_126630_1706# a_126010_2496# a_126520_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X859 word4.byte4.tinv7.O word4.byte4.tinv4.EN a_17220_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X860 a_58050_7978# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X861 VDD word5.byte4.tinv5.I a_20820_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X862 VDD word3.byte1.cgate0.nand0.B word3.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X863 a_93540_12068# word8.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X864 a_121080_7976# buf_out11.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X865 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X866 a_111610_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X867 VDD a_166260_680# a_166220_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X868 word2.byte3.dff_6.O word2.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X869 a_67620_9714# word7.byte3.tinv7.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X870 a_22770_7978# word6.byte4.cgate0.inv1.O a_22660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X871 word3.byte1.tinv7.O buf_out8.inv0.I a_142500_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X872 VSS word3.byte1.cgate0.nand0.B a_73020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X873 a_115440_7978# a_115210_8768# a_114880_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X874 VDD word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X875 a_15460_3326# a_13620_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X876 a_11580_4842# a_11350_5632# a_11020_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X877 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X878 a_154860_6462# word5.byte1.dff_7.CLK a_154300_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X879 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X880 VSS a_155460_680# word1.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X881 VSS word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X882 VDD word3.byte4.tinv5.I a_20820_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X883 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X884 word6.gt_re3.I word6.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X885 a_15780_6952# a_15570_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X886 word5.byte3.cgate0.inv1.I word5.byte3.cgate0.nand0.A a_73020_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X887 a_4770_190# a_4150_140# a_4660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X888 a_11580_1706# a_11350_2496# a_11020_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X889 a_154860_3326# word3.byte1.dff_7.CLK a_154300_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X890 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X891 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X892 VDD word7.byte1.cgate0.nand0.B word7.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X893 a_15780_3816# a_15570_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X894 a_162660_5492# a_162450_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X895 Do22_buf buf_out23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X896 a_15180_10498# a_14950_9548# a_14620_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X897 a_43980_9598# word7.byte3.cgate0.inv1.O a_43420_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X898 a_55340_6462# a_54550_6412# a_55170_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X899 VSS a_8580_2356# word2.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X900 Do3_buf buf_out4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X901 VSS a_162660_11764# word8.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X902 a_7750_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X903 a_6420_4840# word4.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X904 a_166220_7362# word5.byte1.dff_7.CLK a_166050_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X905 a_165660_190# word1.byte1.dff_7.CLK a_165100_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X906 word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.latch0.I0.O a_75720_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X907 a_162340_9048# a_160500_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X908 a_160500_9714# word7.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X909 VSS a_62580_8628# a_62540_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X910 VSS word1.byte4.dff_0.O_bar a_2820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X911 word2.byte1.tinv7.O word2.byte1.tinv5.EN a_160500_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X912 VSS a_147100_11064# a_146100_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X913 a_55340_3326# a_54550_3276# a_55170_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X914 VSS a_114880_7928# a_113880_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X915 a_4940_7978# word6.byte4.cgate0.inv1.O a_4770_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X916 a_108010_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X917 word1.byte1.nand.B word1.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X918 word6.byte4.cgate0.inv1.I word6.byte4.cgate0.nand0.A a_33420_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X919 word1.byte3.tinv7.O word1.byte3.tinv5.EN a_60420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X920 a_166220_4226# word3.byte1.dff_7.CLK a_166050_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X921 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X922 VSS a_57820_1656# a_56820_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X923 a_4660_7362# a_2820_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X924 a_25980_1090# a_25750_140# a_25420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X925 a_147100_7928# word6.byte1.dff_7.CLK a_147330_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X926 VDD word1.byte1.buf_RE1.I word1.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X927 a_108010_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X928 a_105200_4842# word4.byte2.dff_7.CLK a_105030_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X929 VSS buf_sel8.inv0.O buf_sel8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X930 VDD word7.byte2.buf_RE1.I word7.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X931 word5.gt_re3.I word5.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X932 a_113880_6578# word5.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X933 a_4660_4226# a_2820_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X934 word4.byte3.tinv7.O word4.byte3.tinv2.EN a_49620_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X935 VDD buf_ck.inv0.O CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X936 a_105200_1706# word2.byte2.dff_7.CLK a_105030_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X937 word3.gt_re3.I word3.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X938 a_4980_6952# a_4770_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X939 a_140230_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X940 a_153300_7976# buf_out5.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X941 a_53220_6578# word5.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X942 VDD word8.byte3.nand.OUT word8.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X943 word7.byte4.tinv7.O word7.byte4.tinv7.EN a_28020_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X944 buf_out16.inv1.O buf_out16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X945 a_143830_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X946 VSS a_118480_9548# a_117480_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X947 VSS a_14620_6412# a_13620_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X948 a_4980_3816# a_4770_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X949 VSS a_55380_10088# word7.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X950 a_53220_3442# word3.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X951 a_57820_11064# word8.byte3.cgate0.inv1.O a_58050_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X952 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X953 a_146100_9714# buf_out7.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X954 Do27_buf buf_out28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X955 VSS a_10020_4840# a_11580_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X956 VSS a_14620_3276# a_13620_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X957 VSS word6.byte1.tinv1.I a_146100_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X958 VSS a_56820_1704# a_58380_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X959 a_7650_5912# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X960 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X961 a_8540_12184# a_7750_11904# a_8370_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X962 a_119600_1090# word1.byte2.dff_7.CLK a_119430_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X963 VSS buf_out22.inv0.O Do21_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X964 a_141060_8628# a_140850_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X965 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X966 a_40150_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X967 VDD buf_out3.inv0.O Do2_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X968 VSS a_56820_11112# a_58380_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X969 word4.byte1.dff_2.O word4.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X970 VDD a_62580_11764# a_62540_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X971 a_155250_9598# a_154630_9548# a_155140_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X972 VSS word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X973 VSS word3.byte1.cgate0.nand0.B a_134580_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X974 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X975 a_125680_4792# word4.byte2.dff_7.CLK a_125910_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X976 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X977 word2.byte1.dff_2.O word2.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X978 word3.byte1.tinv7.O word3.byte1.tinv1.EN a_146100_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X979 VDD word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X980 VSS a_150700_140# a_149700_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X981 word8.gt_re3.I word8.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X982 VDD buf_we3.inv0.O buf_we3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X983 a_26370_7978# a_25750_8768# a_26260_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X984 a_125680_1656# word2.byte2.dff_7.CLK a_125910_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X985 a_116040_11764# a_115830_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X986 a_155460_10088# a_155250_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X987 VSS word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X988 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X989 VSS a_12180_10088# a_12140_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X990 a_146100_6578# word5.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X991 VDD word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X992 VDD a_3820_6412# a_2820_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X993 buf_in12.inv1.O buf_in12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X994 VSS a_116040_11764# a_116000_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X995 word7.byte3.tinv7.O word7.byte3.tinv5.EN a_60420_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X996 a_64020_4840# buf_out18.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X997 VDD a_121080_9714# a_122640_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X998 a_122410_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X999 VSS a_105240_5492# a_105200_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1000 VDD a_164100_7976# a_165660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1001 a_8370_11114# a_7750_11904# a_8260_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1002 VDD a_15780_10088# word7.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1003 a_151650_9598# word7.byte1.dff_7.CLK a_151540_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1004 VSS word5.byte4.cgate0.nand0.A a_35760_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1005 VDD word6.byte3.tinv6.I a_64020_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1006 VDD a_3820_3276# a_2820_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1007 a_64020_1704# buf_out18.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1008 a_122410_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1009 buf_in6.inv1.O buf_in6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1010 buf_in29.inv1.O buf_in29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1011 a_1380_11764# a_1170_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1012 a_112440_8628# a_112230_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1013 VSS a_1380_6952# a_1340_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1014 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1015 VDD a_66180_8628# a_66140_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1016 a_56820_9714# word7.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1017 VSS word4.byte1.tinv3.I a_153300_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1018 buf_in30.inv1.O buf_in30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1019 VSS buf_in18.inv0.O buf_in18.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1020 VSS a_1380_11764# a_1340_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1021 word8.byte2.tinv7.O buf_out16.inv0.I a_103080_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1022 a_8260_9598# a_6420_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1023 VSS a_100380_190# a_101040_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1024 VSS a_60420_7976# a_61980_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1025 a_122310_190# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1026 VSS a_1380_3816# a_1340_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1027 a_110280_4840# word4.byte2.tinv2.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1028 VDD buf_in21.inv0.O buf_in21.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1029 a_53220_11112# word8.byte3.tinv3.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1030 a_4380_7978# a_4150_8768# a_3820_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1031 word6.byte3.tinv7.O word6.byte3.tinv7.EN a_67620_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1032 a_73020_2660# word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1033 word4.byte3.dff_0.O word4.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1034 word5.byte1.tinv7.O buf_out1.inv0.I a_167700_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1035 VSS buf_sel3.inv0.O buf_sel3.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1036 VDD word5.byte2.tinv3.I a_113880_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1037 a_8580_10088# a_8370_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1038 word1.byte4.tinv7.O buf_out31.inv0.I a_6420_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1039 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1040 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1041 a_70500_13636# dec8.and4_3.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1042 a_147660_9048# word6.byte1.dff_7.CLK a_147100_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1043 a_47970_7978# word6.byte3.cgate0.inv1.O a_47860_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1044 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1045 VSS word7.byte1.nand.B a_39180_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1046 a_140130_9048# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1047 word3.byte1.tinv7.O buf_out1.inv0.I a_167700_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1048 a_18220_4792# a_18550_5632# a_18450_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1049 VDD word3.byte2.tinv3.I a_113880_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1050 VDD a_154300_4792# a_153300_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1051 VDD word4.byte1.cgate0.nand0.A word4.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1052 VDD word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1053 VDD word1.byte3.buf_RE0.O word1.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1054 a_67620_11112# buf_out17.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1055 word6.byte3.dff_5.O word6.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1056 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1057 a_113880_306# word1.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1058 VDD word7.byte1.nand.B word7.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1059 a_56820_3442# word3.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1060 VSS word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1061 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1062 VSS a_107680_140# a_106680_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1063 VDD a_154300_1656# a_153300_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1064 VDD word2.byte1.cgate0.nand0.A word2.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1065 a_13620_3442# word3.byte4.tinv3.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1066 buf_out12.inv1.O buf_out12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1067 VSS a_123240_11764# word8.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1068 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1069 a_48140_9048# a_47350_8768# a_47970_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1070 VSS a_112440_2356# a_112400_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1071 VDD a_19380_11764# a_19340_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1072 VSS a_3820_7928# a_2820_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1073 a_18780_190# word1.byte4.cgate0.inv1.O a_18220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1074 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1075 a_121080_9714# word7.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1076 word1.byte3.dff_2.O word1.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1077 a_14950_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1078 VDD a_43420_7928# a_42420_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1079 a_24420_7976# word6.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1080 a_44260_11114# a_42420_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1081 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1082 a_61650_9598# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1083 VSS word1.buf_ck1.I word1.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1084 a_134580_12068# word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1085 a_118710_7362# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1086 buf_in28.inv1.O buf_in28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1087 VSS word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1088 VSS buf_out3.inv0.I buf_out3.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X1089 word7.byte4.cgate0.nand0.A word7.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1090 a_144660_8628# a_144450_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1091 a_100480_140# word1.byte2.dff_7.CLK a_100710_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1092 VSS a_124680_306# a_126240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1093 VDD a_24420_11112# a_25980_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1094 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1095 a_118710_4226# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1096 Do31_buf buf_out32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1097 VDD buf_out18.inv0.O Do17_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1098 VDD buf_in5.inv0.O buf_in5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1099 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1100 VSS word7.byte1.tinv6.I a_164100_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1101 VDD word7.byte3.tinv5.I a_60420_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1102 VSS buf_we3.inv0.O buf_we3.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1103 a_13620_11112# word8.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1104 a_43650_1090# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1105 a_121080_306# buf_out11.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1106 a_104920_9598# a_103080_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1107 a_140230_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1108 a_111510_7978# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1109 VDD a_48180_5492# word4.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1110 VSS word4.byte3.cgate0.nand0.A a_75360_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1111 VDD buf_sel1.inv0.O buf_sel1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1112 a_148050_11114# a_147430_11904# a_147940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1113 VDD word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1114 VSS a_7420_9548# a_6420_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1115 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1116 VDD a_151860_680# a_151820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1117 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1118 a_154530_12184# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1119 VDD word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1120 a_26370_11114# word8.byte4.cgate0.inv1.O a_26260_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1121 a_101040_7978# a_100810_8768# a_100480_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1122 VDD a_48180_2356# word2.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1123 word1.gt_re3.I word1.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1124 buf_sel5.inv1.O buf_sel5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1125 a_57820_9548# word7.byte3.cgate0.inv1.O a_58050_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1126 a_106680_9714# buf_out15.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1127 word5.byte2.dff_5.O word5.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1128 a_25420_1656# a_25750_2496# a_25650_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1129 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1130 VDD a_7420_11064# a_6420_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1131 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1132 word8.byte3.dff_1.O word8.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1133 VDD word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1134 VSS a_39820_6412# a_39720_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1135 a_220_140# word1.byte4.cgate0.inv1.O a_450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1136 buf_we4.inv1.O buf_we4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1137 a_154300_11064# word8.byte1.dff_7.CLK a_154530_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1138 a_11350_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1139 word3.byte2.dff_5.O word3.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1140 VDD word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1141 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1142 a_44580_11764# a_44370_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1143 a_150700_9548# a_151030_9548# a_150930_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1144 a_105200_190# a_104410_140# a_105030_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1145 buf_re.inv1.O buf_re.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1146 VSS a_39820_3276# a_39720_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1147 a_40940_6462# a_40150_6412# a_40770_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1148 word8.byte1.tinv7.O word8.byte1.tinv1.EN a_146100_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1149 a_11350_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1150 VDD Di24 buf_in25.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1151 VDD buf_out11.inv0.O buf_out11.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1152 a_151820_7362# word5.byte1.dff_7.CLK a_151650_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1153 VDD a_62580_10088# a_62540_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1154 a_128280_8932# word6.byte2.tinv7.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1155 a_134580_2660# word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1156 a_166260_8628# a_166050_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1157 a_40940_3326# a_40150_3276# a_40770_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1158 VSS buf_out2.inv0.O Do1_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1159 a_65350_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1160 a_144450_190# word1.byte1.dff_7.CLK a_144340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1161 a_55380_5492# a_55170_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1162 VSS a_148260_6952# a_148220_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1163 VSS a_153300_11112# a_154860_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1164 VSS word2.gt_re1.O word2.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1165 a_151820_4226# word3.byte1.dff_7.CLK a_151650_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1166 Do30_buf buf_out31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1167 word1.byte4.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1168 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1169 a_116040_10088# a_115830_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1170 a_55380_2356# a_55170_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1171 VSS a_148260_3816# a_148220_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1172 a_144450_4842# a_143830_5632# a_144340_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1173 VDD a_112440_8628# word6.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1174 a_53220_1704# word2.byte3.tinv3.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1175 VSS word3.byte2.tinv4.I a_117480_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1176 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1177 a_119430_1706# word2.byte2.dff_7.CLK a_119320_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1178 Do16_buf buf_out17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1179 a_153300_306# buf_out5.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1180 word3.byte1.nand.OUT buf_we4.inv1.O a_129540_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1181 a_8370_9598# a_7750_9548# a_8260_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1182 a_144450_1706# a_143830_2496# a_144340_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1183 VSS word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1184 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1185 word3.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1186 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1187 VSS word3.byte1.cgate0.nand0.B word3.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1188 VDD word6.byte1.buf_RE1.I word6.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1189 VDD word5.byte4.nand.OUT word5.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1190 VSS a_20820_306# a_22380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1191 a_35760_4840# word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1192 a_1380_10088# a_1170_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1193 VSS word3.byte4.inv_and.O a_36120_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1194 buf_in14.inv1.O buf_in14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1195 VSS a_40980_10088# word7.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1196 word6.byte1.nand.B word6.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1197 a_35760_1704# word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1198 VDD word3.byte4.nand.OUT word3.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1199 VDD word7.byte4.tinv4.I a_17220_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1200 buf_in28.inv1.O buf_in28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1201 VDD a_19380_680# a_19340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1202 a_61420_6412# a_61750_6412# a_61650_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1203 VSS word6.byte1.inv_and.O a_131700_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1204 a_15460_5912# a_13620_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1205 VSS word8.byte2.tinv6.I a_124680_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1206 word7.byte3.tinv7.O buf_out24.inv0.I a_42420_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1207 a_62260_190# a_60420_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1208 a_61420_3276# a_61750_3276# a_61650_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1209 a_158850_190# a_158230_140# a_158740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1210 VSS buf_in20.inv0.O buf_in20.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1211 VDD a_22980_680# word1.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1212 word6.byte2.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B a_93540_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1213 a_20820_306# word1.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1214 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1215 a_154860_5912# word4.byte1.dff_7.CLK a_154300_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1216 VSS word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1217 a_149700_11112# word8.byte1.tinv2.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1218 a_2820_9714# word7.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1219 VDD buf_we2.inv0.O buf_we2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1220 a_39180_8932# buf_we1.inv1.O word6.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1221 a_15780_5492# a_15570_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1222 word2.byte2.dff_2.O word2.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1223 a_111280_4792# word4.byte2.dff_7.CLK a_111510_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1224 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1225 a_75720_10500# word7.byte3.cgate0.latch0.I0.ENB word7.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1226 VDD word5.byte1.buf_RE1.I word5.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1227 VSS dec8.and4_5.nand0.OUT buf_sel6.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1228 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1229 VDD EN dec8.and4_5.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1230 a_19340_7362# word5.byte4.cgate0.inv1.O a_19170_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1231 VDD word4.byte1.tinv5.I a_160500_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1232 VDD buf_sel8.inv0.O buf_sel8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1233 VSS word8.buf_sel0.O word8.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1234 a_11970_7978# a_11350_8768# a_11860_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1235 a_6420_6578# word5.byte4.tinv1.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1236 VSS word7.byte3.inv_and.O a_75720_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1237 a_165330_9048# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1238 a_111280_1656# word2.byte2.dff_7.CLK a_111510_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1239 word2.byte4.tinv7.O word2.byte4.tinv3.EN a_13620_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1240 VDD word3.byte1.buf_RE1.I word3.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1241 a_55340_5912# a_54550_5632# a_55170_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1242 a_164100_11112# buf_out2.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1243 a_54450_4842# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1244 a_131700_6578# word5.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1245 word6.byte4.dff_6.O word6.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1246 VDD a_149700_306# a_151260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1247 a_158230_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1248 VDD a_19380_10088# a_19340_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1249 VDD word2.byte1.tinv5.I a_160500_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1250 VSS a_46020_306# a_47580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1251 a_19340_4226# word3.byte4.cgate0.inv1.O a_19170_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1252 VDD word4.byte1.nand.OUT word4.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1253 word4.byte2.tinv7.O buf_out12.inv0.I a_117480_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1254 a_158740_7362# a_156900_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1255 VDD a_58980_6952# a_58940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1256 VSS word5.buf_ck1.I word5.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1257 VDD word1.byte3.tinv6.I a_64020_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1258 VDD a_162660_5492# a_162620_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1259 a_44260_10498# a_42420_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1260 a_54450_190# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1261 a_54450_1706# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1262 a_93540_6578# word5.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1263 a_108010_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1264 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1265 a_12140_7978# word6.byte4.cgate0.inv1.O a_11970_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1266 a_160500_306# word1.byte1.tinv5.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1267 a_10020_7976# word6.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1268 a_147430_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1269 VDD word2.byte1.nand.OUT word2.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1270 word2.byte2.tinv7.O buf_out12.inv0.I a_117480_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1271 a_158740_4226# a_156900_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1272 VSS buf_out11.inv0.I buf_out11.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X1273 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1274 a_155420_9598# a_154630_9548# a_155250_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1275 VDD a_162660_2356# a_162620_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1276 VDD a_58980_3816# a_58940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1277 a_49620_7976# word6.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1278 a_61650_11114# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1279 a_115440_12184# word8.byte2.dff_7.CLK a_114880_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1280 VDD a_24420_9714# a_25980_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1281 VSS a_108840_8628# a_108800_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1282 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1283 Do6_buf buf_out7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1284 a_126800_11114# word8.byte2.dff_7.CLK a_126630_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1285 a_151540_7978# a_149700_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1286 a_40380_6462# word5.byte3.cgate0.inv1.O a_39820_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1287 a_44580_680# a_44370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1288 a_106680_306# word1.byte2.tinv1.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1289 VDD a_51780_8628# a_51740_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1290 a_164100_7976# word6.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1291 Do30_buf buf_out31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1292 VSS buf_in4.inv0.O buf_in4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1293 a_4150_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1294 a_22660_2776# a_20820_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1295 a_151260_7362# a_151030_6412# a_150700_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1296 a_51570_6462# a_50950_6412# a_51460_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1297 a_46020_306# word1.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1298 VSS a_157900_4792# a_156900_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1299 VSS word4.byte1.buf_RE1.I word4.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1300 a_40380_3326# word3.byte3.cgate0.inv1.O a_39820_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1301 VDD buf_out22.inv0.I buf_out22.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X1302 a_108630_11114# a_108010_11904# a_108520_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1303 a_148050_9598# a_147430_9548# a_147940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1304 word5.byte3.dff_6.O word5.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1305 word6.byte3.tinv7.O word6.byte3.tinv3.EN a_53220_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1306 a_1340_4842# word4.byte4.cgate0.inv1.O a_1170_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1307 a_4150_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1308 a_115110_12184# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1309 a_151260_4226# a_151030_3276# a_150700_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1310 a_51570_3326# a_50950_3276# a_51460_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1311 word5.byte1.tinv7.O buf_out5.inv0.I a_153300_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1312 VDD word8.byte1.cgate0.nand0.A word8.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1313 a_7980_12184# word8.byte4.cgate0.inv1.O a_7420_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1314 word1.byte3.cgate0.nand0.A word1.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1315 a_22980_2356# a_22770_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1316 word3.byte3.dff_6.O word3.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1317 a_12140_190# a_11350_140# a_11970_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1318 a_126240_1090# a_126010_140# a_125680_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1319 a_1340_1706# word2.byte4.cgate0.inv1.O a_1170_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1320 a_60420_11112# word8.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1321 VDD word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1322 word7.byte3.dff_1.O word7.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1323 word6.byte2.dff_3.O word6.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1324 VSS a_166260_8628# word6.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1325 word3.byte1.tinv7.O buf_out5.inv0.I a_153300_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1326 a_110280_3442# word3.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1327 a_114880_11064# word8.byte2.dff_7.CLK a_115110_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1328 a_154300_9548# word7.byte1.dff_7.CLK a_154530_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1329 a_36120_9714# word7.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1330 VSS a_108840_11764# a_108800_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1331 VSS word5.gt_re1.O word5.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1332 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1333 a_62540_2776# a_61750_2496# a_62370_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1334 word8.byte1.dff_7.O word8.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1335 VDD a_8580_6952# word5.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1336 word8.byte2.tinv7.O word8.byte2.tinv1.EN a_106680_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1337 VSS word5.byte4.buf_RE0.O word5.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1338 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1339 word4.gt_re1.O word4.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1340 a_24420_306# word1.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1341 a_140230_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1342 a_141060_11764# a_140850_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1343 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1344 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1345 VDD word4.byte4.tinv7.I a_28020_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1346 a_115210_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1347 VDD a_8580_3816# word3.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1348 VDD a_148260_11764# word8.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1349 VDD a_154300_9548# a_153300_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1350 word2.gt_re1.O word2.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1351 buf_in10.inv0.O buf_in10.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1352 a_140230_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1353 buf_we1.inv1.O buf_we1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1354 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B a_132960_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1355 VDD word2.byte4.tinv7.I a_28020_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1356 buf_in1.inv0.O Di0 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1357 VDD a_1380_8628# word6.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1358 VSS buf_we2.inv0.O buf_we2.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1359 VDD a_17220_7976# a_18780_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1360 a_118810_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1361 a_117480_1704# word2.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1362 a_8370_1706# word2.byte4.cgate0.inv1.O a_8260_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1363 buf_in30.inv1.O buf_in30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1364 a_46020_11112# word8.byte3.tinv1.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1365 a_157900_140# word1.byte1.dff_7.CLK a_158130_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1366 VDD buf_out27.inv0.I buf_out27.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X1367 a_129540_2660# word2.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1368 VDD a_11020_6412# a_10020_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1369 a_118810_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1370 a_116000_4842# word4.byte2.dff_7.CLK a_115830_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1371 a_149700_9714# word7.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1372 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1373 VDD a_11020_3276# a_10020_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1374 a_18450_11114# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1375 VSS word7.byte2.buf_RE1.I word7.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1376 word7.byte2.tinv7.O word7.byte2.tinv1.EN a_106680_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1377 a_116000_1706# word2.byte2.dff_7.CLK a_115830_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1378 word1.byte2.dff_6.O word1.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1379 a_164100_7976# buf_out2.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1380 a_64020_6578# word5.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1381 a_154630_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1382 VSS a_1380_5492# a_1340_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1383 a_20820_6578# buf_out27.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1384 VSS a_116040_11764# word8.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1385 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1386 VSS word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1387 a_64020_3442# word3.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1388 VDD a_56820_6578# a_58380_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1389 VDD word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1390 a_54220_7928# a_54550_8768# a_54450_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1391 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1392 VDD a_160500_4840# a_162060_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1393 a_113880_9714# word7.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1394 VSS a_162660_680# word1.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1395 VSS buf_in13.inv0.O buf_in13.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1396 word8.byte3.inv_and.O word8.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1397 VSS word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1398 a_20820_3442# buf_out27.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1399 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1400 VDD word6.byte4.buf_RE0.O word6.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1401 VDD word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1402 VDD a_56820_3442# a_58380_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1403 a_110280_11112# word8.byte2.tinv2.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1404 a_55170_9598# word7.byte3.cgate0.inv1.O a_55060_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1405 VDD a_160500_1704# a_162060_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1406 a_17220_11112# word8.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1407 word1.byte1.nand.OUT buf_we4.inv1.O a_129540_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1408 a_25650_6462# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1409 a_113880_7976# word6.byte2.tinv3.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1410 VSS a_108840_680# word1.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1411 word7.byte3.dff_7.O word7.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1412 VDD a_17220_11112# a_18780_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1413 a_50950_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1414 VDD a_49620_7976# a_51180_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1415 VDD a_107680_11064# a_106680_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1416 a_25650_3326# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1417 VDD buf_in24.inv0.O buf_in24.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1418 word4.byte4.tinv7.O word4.byte4.tinv1.EN a_6420_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1419 a_75720_8932# word6.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1420 VSS word2.byte3.buf_RE0.O word2.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1421 a_82020_2660# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1422 a_55340_12184# a_54550_11904# a_55170_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1423 a_76620_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1424 a_124680_11112# buf_out10.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1425 VSS a_121080_6578# a_122640_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1426 a_158230_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1427 VSS word6.byte1.cgate0.nand0.B a_33420_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1428 VSS word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1429 VSS word4.byte3.buf_RE0.O word4.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1430 a_105030_1706# word2.byte2.dff_7.CLK a_104920_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1431 a_148220_4842# word4.byte1.dff_7.CLK a_148050_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1432 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1433 word1.byte3.dff_2.O word1.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1434 VSS a_11020_7928# a_10020_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1435 word6.byte2.dff_4.O word6.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1436 VSS a_22980_10088# a_22940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1437 VDD word1.byte1.buf_RE1.I word1.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1438 VSS a_121080_3442# a_122640_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1439 a_156900_6578# word5.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1440 a_104640_190# word1.byte2.dff_7.CLK a_104080_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1441 word5.gt_re3.I word5.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1442 VSS word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1443 a_13620_306# word1.byte4.tinv3.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1444 a_148220_1706# word2.byte1.dff_7.CLK a_148050_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1445 word5.byte2.tinv7.O word5.byte2.tinv3.EN a_113880_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1446 word1.byte1.nand.B word1.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1447 a_61650_10498# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1448 VSS word7.byte4.tinv4.I a_17220_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1449 buf_out15.inv1.O buf_out15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1450 word3.gt_re3.I word3.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1451 a_126800_10498# word7.byte2.dff_7.CLK a_126630_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1452 a_4150_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1453 a_107910_9598# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1454 Do5_buf buf_out6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1455 a_123240_680# a_123030_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1456 VDD word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1457 a_55170_11114# a_54550_11904# a_55060_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1458 a_33420_6578# word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1459 word8.byte2.inv_and.O word8.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1460 a_108630_9598# a_108010_9548# a_108520_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1461 a_65580_6462# word5.byte3.cgate0.inv1.O a_65020_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1462 a_47860_2776# a_46020_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1463 a_65580_3326# word3.byte3.cgate0.inv1.O a_65020_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1464 a_121080_4840# word4.byte2.tinv5.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1465 word4.byte2.dff_5.O word4.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1466 VSS word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1467 VDD word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1468 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1469 VSS a_39820_4792# a_39720_4842# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1470 buf_in18.inv1.O buf_in18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1471 a_114880_9548# word7.byte2.dff_7.CLK a_115110_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1472 VDD word5.byte2.tinv6.I a_124680_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1473 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1474 a_93540_306# word1.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1475 a_48180_2356# a_47970_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1476 word4.gt_re3.I word4.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1477 word7.byte1.inv_and.O word7.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1478 word8.byte2.dff_0.O word8.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1479 a_101320_6462# a_100380_6462# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1480 word7.byte1.dff_7.O word7.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1481 a_150930_9048# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1482 a_19380_8628# a_19170_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1483 VDD word3.byte2.tinv6.I a_124680_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1484 a_40940_5912# a_40150_5632# a_40770_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1485 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1486 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1487 CLK buf_ck.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1488 a_101640_11764# a_101430_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1489 VDD a_112440_6952# a_112400_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1490 VSS a_139900_9548# a_139800_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1491 a_101320_3326# a_100380_3326# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1492 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1493 word4.byte2.tinv7.O buf_out16.inv0.I a_103080_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1494 VDD word4.byte2.cgate0.nand0.A word4.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1495 a_95160_12068# word8.byte2.cgate0.nand0.A word8.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1496 VDD a_148260_10088# word7.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1497 VSS word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1498 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1499 VSS a_120_6462# a_780_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1500 a_49620_306# word1.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1501 a_57820_7928# word6.byte3.cgate0.inv1.O a_58050_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1502 VDD a_112440_3816# a_112400_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1503 a_165430_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1504 VSS a_148260_5492# a_148220_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1505 word8.byte3.tinv7.O buf_out19.inv0.I a_60420_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1506 a_58940_9048# a_58150_8768# a_58770_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1507 word6.byte2.cgate0.inv1.I word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1508 a_103080_7976# word6.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1509 word2.byte2.tinv7.O buf_out16.inv0.I a_103080_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1510 VDD word2.byte2.cgate0.nand0.A word2.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1511 VSS a_108840_10088# word7.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1512 a_141020_9598# a_140230_9548# a_140850_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1513 buf_in9.inv0.O buf_in9.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1514 VSS word5.byte4.tinv6.I a_24420_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1515 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1516 VSS a_120_3326# a_780_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1517 a_165430_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1518 VDD buf_out14.inv0.O buf_out14.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1519 VSS word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1520 VDD word7.byte4.cgate0.nand0.A a_35760_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1521 a_155460_8628# a_155250_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1522 VSS buf_out5.inv0.O Do4_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1523 a_54550_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1524 VDD buf_in5.inv0.O buf_in5.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1525 VSS a_66180_680# a_66140_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1526 a_167700_12068# word8.byte1.tinv7.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1527 buf_in20.inv0.O Di19 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1528 a_18450_10498# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1529 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1530 a_122310_1090# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1531 a_51460_9048# a_49620_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1532 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1533 a_153300_4840# word4.byte1.tinv3.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1534 VSS dec8.and4_1.nand0.OUT buf_sel2.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1535 VDD a_58980_5492# word4.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1536 a_111840_1090# a_111610_140# a_111280_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1537 a_25420_6412# word5.byte4.cgate0.inv1.O a_25650_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1538 VSS a_62580_11764# word8.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1539 VDD word5.byte1.tinv4.I a_156900_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1540 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1541 VSS a_151860_8628# word6.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1542 VDD a_58980_2356# word2.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1543 VDD word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1544 a_61420_4792# a_61750_5632# a_61650_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1545 VSS buf_sel6.inv0.I buf_sel6.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1546 a_51780_8628# a_51570_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1547 word5.byte4.cgate0.nand0.A word5.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1548 a_147940_190# a_146100_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1549 a_104080_1656# a_104410_2496# a_104310_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1550 VSS word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1551 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1552 a_25420_3276# word3.byte4.cgate0.inv1.O a_25650_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1553 VSS a_20820_9714# a_22380_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1554 VDD word3.byte1.tinv4.I a_156900_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1555 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1556 a_22150_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1557 a_46020_6578# buf_out23.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1558 buf_sel1.inv1.O buf_sel1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1559 a_119640_680# a_119430_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1560 VSS word3.byte2.buf_RE1.I word3.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1561 word3.byte4.cgate0.nand0.A word3.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1562 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1563 a_47250_2776# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1564 VDD word7.byte2.buf_RE1.I word7.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1565 a_161500_9548# a_161830_9548# a_161730_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1566 VSS a_100480_6412# a_100380_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1567 word3.byte3.tinv7.O word3.byte3.tinv4.EN a_56820_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1568 a_46020_3442# buf_out23.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1569 VDD word4.byte4.tinv3.I a_13620_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1570 a_151540_11114# a_149700_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1571 VDD a_54220_11064# a_53220_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1572 VDD a_17220_9714# a_18780_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1573 a_18450_9048# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1574 VSS a_155460_2356# a_155420_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1575 a_100810_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1576 VSS a_114880_140# a_113880_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1577 VDD buf_in10.inv0.O buf_in10.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1578 VSS a_100480_3276# a_100380_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1579 VDD a_154300_140# a_153300_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1580 VDD word2.byte4.tinv3.I a_13620_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1581 a_25980_190# word1.byte4.cgate0.inv1.O a_25420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1582 word1.byte3.dff_4.O word1.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1583 VSS buf_in29.inv0.O buf_in29.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1584 VSS a_4980_680# a_4940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1585 VSS buf_in23.inv0.O buf_in23.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1586 VDD buf_we1.inv1.O word7.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1587 word6.byte4.tinv7.O buf_out26.inv0.I a_24420_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1588 a_108240_6462# word5.byte2.dff_7.CLK a_107680_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1589 VDD a_15780_5492# a_15740_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1590 VDD buf_in4.inv0.O buf_in4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1591 a_119430_6462# a_118810_6412# a_119320_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1592 a_143500_140# word1.byte1.dff_7.CLK a_143730_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1593 VSS a_113880_7976# a_115440_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1594 word2.byte4.dff_1.O word2.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1595 a_107910_12184# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1596 a_151820_12184# a_151030_11904# a_151650_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1597 VDD a_123240_680# word1.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1598 VDD a_15780_2356# a_15740_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1599 a_108240_3326# word3.byte2.dff_7.CLK a_107680_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1600 a_64020_1704# word2.byte3.tinv6.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1601 a_119430_3326# a_118810_3276# a_119320_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1602 VSS a_116040_10088# a_116000_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1603 a_164100_306# buf_out2.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1604 a_147940_9598# a_146100_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1605 a_154530_7978# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1606 word2.byte1.dff_5.O word2.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1607 a_17220_7976# word6.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1608 VSS word4.byte3.tinv6.I a_64020_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1609 VDD word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1610 buf_sel4.inv0.I dec8.and4_3.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1611 a_4150_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1612 a_112230_7978# a_111610_8768# a_112120_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1613 a_40380_5912# word4.byte3.cgate0.inv1.O a_39820_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1614 VDD buf_sel7.inv0.I buf_sel7.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1615 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1616 word4.byte4.dff_5.O word4.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1617 a_4150_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1618 buf_in14.inv1.O buf_in14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1619 a_55170_9598# a_54550_9548# a_55060_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1620 word5.byte1.dff_6.O word5.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1621 VSS word5.buf_sel0.O word5.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1622 a_159060_11764# a_158850_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1623 VDD word1.byte4.buf_RE0.O word1.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1624 a_139900_11064# a_140230_11904# a_140130_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1625 VSS a_4980_8628# a_4940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1626 word2.byte4.dff_5.O word2.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1627 VSS buf_out12.inv0.O buf_out12.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1628 VDD a_100480_11064# a_100380_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1629 a_58380_9048# word6.byte3.cgate0.inv1.O a_57820_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1630 word3.byte1.dff_6.O word3.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1631 VSS a_124680_11112# a_126240_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1632 a_140460_9598# word7.byte1.dff_7.CLK a_139900_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1633 a_40770_9598# word7.byte3.cgate0.inv1.O a_40660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1634 VDD a_65020_4792# a_64020_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1635 VDD word8.gt_re1.O word8.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1636 a_112400_190# a_111610_140# a_112230_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1637 word7.byte3.dff_3.O word7.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1638 word5.byte2.dff_2.O word5.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1639 VDD a_65020_1656# a_64020_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1640 VDD buf_out1.inv0.O Do0_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1641 VDD buf_out23.inv0.O Do22_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1642 word7.byte2.dff_0.O word7.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1643 a_55060_7978# a_53220_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1644 VSS a_154300_1656# a_153300_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1645 a_134580_2660# word2.byte1.cgate0.nand0.A word2.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1646 word3.byte2.dff_2.O word3.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1647 VSS word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1648 VSS buf_out32.inv0.O Do31_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1649 a_22770_190# a_22150_140# a_22660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1650 a_151650_190# word1.byte1.dff_7.CLK a_151540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1651 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1652 a_65100_13636# dec8.and4_0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1653 a_126520_6462# a_124680_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1654 word6.byte2.dff_0.O word6.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1655 VDD a_155460_8628# word6.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1656 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1657 VDD word8.byte1.inv_and.O a_131700_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1658 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1659 a_108800_2776# a_108010_2496# a_108630_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1660 buf_sel1.inv1.O buf_sel1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1661 VDD word8.byte1.cgate0.nand0.B word8.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1662 VDD word8.byte1.tinv4.I a_156900_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1663 VSS a_26580_2356# word2.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1664 a_25750_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1665 a_117480_3442# word3.byte2.tinv4.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1666 word4.byte2.tinv7.O buf_out9.inv0.I a_128280_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1667 VSS a_43420_4792# a_42420_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1668 a_126520_3326# a_124680_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1669 a_122640_4842# a_122410_5632# a_122080_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1670 a_24420_4840# word4.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1671 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1672 word8.gt_re0.OUT buf_sel8.inv1.O a_82020_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1673 a_73020_306# word1.byte3.cgate0.nand0.A word1.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1674 a_118810_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1675 VDD buf_we2.inv1.O word4.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1676 VSS word3.buf_ck1.I word3.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1677 VDD word4.byte2.nand.OUT word4.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1678 a_22940_7978# word6.byte4.cgate0.inv1.O a_22770_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1679 a_128280_7976# word6.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1680 VDD word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1681 word2.byte2.tinv7.O buf_out9.inv0.I a_128280_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1682 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1683 a_122640_1706# a_122410_2496# a_122080_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1684 VSS word5.byte3.tinv2.I a_49620_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1685 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1686 VSS buf_we4.inv0.O buf_we4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1687 a_36120_4840# word4.byte4.cgate0.latch0.I0.ENB word4.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1688 a_22660_7362# a_20820_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1689 a_162340_1090# a_160500_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1690 word6.byte3.inv_and.O word6.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1691 word6.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1692 VDD a_62580_680# a_62540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1693 VDD buf_we2.inv1.O word2.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1694 VDD word2.byte2.nand.OUT word2.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1695 VDD buf_in13.inv0.O buf_in13.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1696 a_103080_11112# word8.byte2.tinv0.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1697 a_128280_12068# word8.byte2.tinv7.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1698 VDD word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1699 a_19170_6462# word5.byte4.cgate0.inv1.O a_19060_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1700 a_36120_1704# word2.byte4.cgate0.latch0.I0.ENB word2.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1701 word7.byte1.tinv7.O buf_out4.inv0.I a_156900_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1702 a_22660_4226# a_20820_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1703 VSS buf_in4.inv0.O buf_in4.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1704 VDD word7.byte4.buf_RE0.O word7.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1705 a_131700_8932# word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1706 a_22980_6952# a_22770_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1707 VDD buf_out30.inv0.O Do29_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1708 VDD a_117480_7976# a_119040_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1709 a_19170_3326# word3.byte4.cgate0.inv1.O a_19060_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1710 VDD a_13620_4840# a_15180_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1711 VSS word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1712 VSS a_156900_6578# a_158460_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1713 a_101640_2356# a_101430_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1714 Do18_buf buf_out19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1715 word6.byte2.cgate0.nand0.A word6.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1716 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1717 a_22980_3816# a_22770_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1718 VDD a_13620_1704# a_15180_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1719 word7.byte4.tinv7.O word7.byte4.tinv0.EN a_2820_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1720 VSS a_156900_3442# a_158460_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1721 a_154300_4792# word4.byte1.dff_7.CLK a_154530_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1722 dec8.and4_7.nand1.OUT A2 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1723 a_62540_7362# word5.byte3.cgate0.inv1.O a_62370_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1724 VSS buf_out17.inv0.O Do16_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1725 a_105240_6952# a_105030_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1726 VSS buf_sel3.inv0.I buf_sel3.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1727 VSS a_46020_9714# a_47580_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1728 VDD word6.byte4.tinv1.I a_6420_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1729 a_154300_1656# word2.byte1.dff_7.CLK a_154530_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1730 a_54780_12184# word8.byte3.cgate0.inv1.O a_54220_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1731 VSS word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1732 a_62540_4226# word3.byte3.cgate0.inv1.O a_62370_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1733 a_151540_10498# a_149700_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1734 a_160500_4840# buf_out3.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1735 a_25650_5912# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1736 word8.byte2.cgate0.nand0.A word8.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1737 a_112120_11114# a_110280_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1738 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1739 a_115210_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1740 word1.byte2.cgate0.inv1.I word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1741 a_103080_306# word1.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1742 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1743 VSS word7.byte1.cgate0.nand0.B word7.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1744 a_112400_9048# a_111610_8768# a_112230_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1745 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1746 a_105240_3816# a_105030_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1747 VSS word3.gt_re0.OUT word3.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1748 VDD word5.byte4.buf_RE0.O word5.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1749 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.latch0.I0.O a_131700_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1750 a_43420_7928# word6.byte3.cgate0.inv1.O a_43650_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1751 VDD word6.buf_ck1.I word6.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1752 VSS buf_in16.inv0.O buf_in16.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1753 VDD a_8580_8628# a_8540_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1754 VSS a_125680_6412# a_124680_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1755 a_160500_1704# buf_out3.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1756 VSS a_62580_6952# word5.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1757 VSS a_53220_306# a_54780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1758 a_115210_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1759 VDD a_150700_11064# a_149700_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1760 word5.gt_re0.OUT buf_sel5.inv1.O a_82020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1761 a_47970_11114# a_47350_11904# a_47860_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1762 a_8370_6462# a_7750_6412# a_8260_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1763 VDD word3.byte4.buf_RE0.O word3.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1764 a_61650_190# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1765 VSS a_121080_4840# a_122640_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1766 VSS a_2820_7976# a_4380_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1767 a_141060_680# a_140850_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1768 VSS a_125680_3276# a_124680_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1769 a_780_4842# a_550_5632# a_220_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1770 a_49620_7976# buf_out22.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1771 a_40150_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1772 a_154630_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1773 VSS a_62580_3816# word3.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1774 a_112400_12184# a_111610_11904# a_112230_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1775 VSS buf_out23.inv0.I buf_out23.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X1776 a_8370_3326# a_7750_3276# a_8260_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1777 a_4660_11114# a_2820_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1778 VDD buf_in26.inv0.O buf_in26.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1779 VSS word8.byte4.tinv3.I a_13620_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1780 a_66180_11764# a_65970_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1781 a_780_1706# a_550_2496# a_220_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1782 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1783 VDD a_21820_6412# a_20820_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1784 a_51780_680# a_51570_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1785 a_113880_306# word1.byte2.tinv3.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1786 VSS a_40980_11764# a_40940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1787 a_160500_9714# buf_out3.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1788 a_1170_7978# a_550_8768# a_1060_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1789 buf_we2.inv1.O buf_we2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1790 VSS a_66180_11764# a_66140_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1791 VSS word6.byte3.dff_0.O_bar a_42420_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1792 a_35760_2660# word2.byte1.cgate0.nand0.B word2.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1793 VSS word4.byte1.buf_RE1.I word4.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1794 VDD a_21820_3276# a_20820_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1795 VDD buf_in32.inv0.O buf_in32.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1796 buf_in18.inv1.O buf_in18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1797 VDD word5.byte1.tinv0.I a_142500_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1798 word4.byte1.nand.B word4.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1799 buf_sel8.inv1.O buf_sel8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1800 VDD word5.byte2.inv_and.O a_92280_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1801 VSS word1.byte1.tinv4.I a_156900_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1802 word6.byte1.dff_4.O word6.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1803 a_65580_5912# word4.byte3.cgate0.inv1.O a_65020_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1804 a_153300_3442# word3.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1805 VDD word3.byte1.tinv0.I a_142500_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1806 word4.byte3.dff_1.O word4.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1807 VDD buf_ck.inv0.I buf_ck.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1808 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1809 VDD a_100480_9548# a_100380_9598# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1810 a_26260_9598# a_24420_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1811 a_4050_9598# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1812 VSS word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1813 VDD word3.byte2.inv_and.O a_92280_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1814 word8.byte3.tinv7.O buf_out21.inv0.I a_53220_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1815 word7.byte4.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1816 word2.byte3.dff_1.O word2.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1817 a_22380_7978# a_22150_8768# a_21820_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1818 word8.byte4.dff_1.O word8.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1819 a_165660_9598# word7.byte1.dff_7.CLK a_165100_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1820 a_104310_6462# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1821 VDD buf_out16.inv0.O buf_out16.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1822 a_65970_9598# word7.byte3.cgate0.inv1.O a_65860_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1823 VSS a_220_1656# a_120_1706# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1824 VDD buf_out9.inv0.O buf_out9.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1825 a_42420_6578# word5.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1826 word1.byte4.tinv7.O buf_out26.inv0.I a_24420_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1827 a_158230_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1828 a_26580_10088# a_26370_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1829 VDD a_60420_306# a_61980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1830 a_4980_11764# a_4770_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1831 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1832 VSS buf_out7.inv0.O Do6_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1833 a_101320_5912# a_100380_4842# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1834 VSS buf_out28.inv0.I buf_out28.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X1835 word6.byte4.tinv7.O buf_out30.inv0.I a_10020_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1836 a_104310_3326# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1837 VSS word2.byte1.tinv5.I a_160500_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1838 a_18550_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1839 a_15740_11114# word8.byte4.cgate0.inv1.O a_15570_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1840 a_105030_6462# a_104410_6412# a_104920_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1841 a_66140_9598# a_65350_9548# a_65970_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1842 a_147660_1090# a_147430_140# a_147100_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1843 a_119320_9048# a_117480_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1844 a_47970_190# a_47350_140# a_47860_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1845 VSS a_120_4842# a_780_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1846 a_140130_1090# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1847 word2.byte2.tinv7.O word2.byte2.tinv4.EN a_117480_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1848 a_18550_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1849 VSS word2.byte1.nand.OUT word2.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1850 a_105030_3326# a_104410_3276# a_104920_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1851 a_159020_4842# word4.byte1.dff_7.CLK a_158850_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1852 buf_in2.inv1.O buf_in2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1853 VSS a_101640_10088# a_101600_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1854 word1.byte3.dff_5.O word1.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1855 VDD EN dec8.and4_2.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1856 word6.byte2.dff_7.O word6.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1857 VSS a_21820_7928# a_20820_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1858 a_149700_9714# word7.byte1.tinv2.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1859 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1860 VDD word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1861 a_22380_11114# a_22150_11904# a_21820_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1862 a_159020_1706# word2.byte1.dff_7.CLK a_158850_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1863 a_49620_4840# word4.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1864 a_14950_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1865 a_44540_190# a_43750_140# a_44370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1866 a_48140_1090# word1.byte3.cgate0.inv1.O a_47970_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1867 word5.byte3.tinv7.O buf_out18.inv0.I a_64020_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1868 VSS buf_in12.inv0.O buf_in12.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1869 word7.byte2.tinv7.O buf_out12.inv0.I a_117480_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1870 VDD word4.byte1.cgate0.nand0.B word4.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1871 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1872 a_47860_7362# a_46020_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1873 a_43980_9048# word6.byte3.cgate0.inv1.O a_43420_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1874 VSS word1.byte4.nand.OUT word1.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1875 a_22660_12184# a_20820_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1876 a_7750_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1877 VDD a_6420_7976# a_7980_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1878 VSS a_105240_6952# word5.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1879 word3.byte3.tinv7.O buf_out18.inv0.I a_64020_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1880 VDD a_50620_4792# a_49620_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1881 VDD word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1882 buf_in32.inv1.O buf_in32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1883 word6.byte3.cgate0.inv1.I word6.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1884 VDD word2.byte1.cgate0.nand0.B word2.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1885 a_47860_4226# a_46020_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1886 VSS buf_we1.inv0.O buf_we1.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1887 VSS buf_in10.inv0.I buf_in10.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1888 VSS a_25420_9548# a_24420_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1889 a_156900_7976# word6.byte1.tinv4.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1890 VSS a_105240_3816# word3.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1891 a_48180_6952# a_47970_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1892 VDD a_50620_1656# a_49620_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X1893 VDD word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1894 a_151860_5492# a_151650_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1895 buf_in29.inv0.O Di28 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1896 VSS a_47020_140# a_46020_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X1897 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1898 a_40660_7978# a_39720_7978# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1899 a_14620_9548# a_14950_9548# a_14850_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1900 a_780_190# word1.byte4.cgate0.inv1.O a_220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1901 word7.byte4.tinv7.O buf_out32.inv0.I a_2820_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1902 VSS a_116040_680# word1.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1903 a_126840_2356# a_126630_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1904 a_56820_9714# buf_out20.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1905 VSS buf_in30.inv0.O buf_in30.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1906 buf_in18.inv1.O buf_in18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1907 a_48180_3816# a_47970_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1908 a_151860_2356# a_151650_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1909 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1910 a_112120_10498# a_110280_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1911 VSS a_100480_4792# a_100380_4842# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1912 VDD Di20 buf_in21.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1913 word6.byte3.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1914 VDD a_141060_8628# word6.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1915 word2.gt_re1.O word2.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1916 VDD word8.byte1.nand.OUT word8.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1917 a_40980_8628# a_40770_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1918 a_148050_1706# word2.byte1.dff_7.CLK a_147940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1919 buf_sel4.inv1.O buf_sel4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1920 VSS word2.byte4.tinv7.I a_28020_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1921 a_103080_3442# word3.byte2.tinv0.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1922 word5.byte1.cgate0.inv1.I word5.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1923 a_128280_1092# word1.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1924 dec8.and4_4.nand0.OUT dec8.and4_6.nand0.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1925 a_47970_9598# a_47350_9548# a_47860_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1926 a_108240_5912# word4.byte2.dff_7.CLK a_107680_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1927 word8.byte4.dff_6.O word8.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1928 VSS word7.byte3.tinv5.I a_60420_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1929 VSS a_55380_8628# word6.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1930 word5.byte1.tinv7.O word5.byte1.tinv4.EN a_156900_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1931 word8.byte3.dff_2.O word8.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1932 VSS word5.byte2.tinv0.I a_103080_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1933 a_113880_7976# word6.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1934 word1.byte3.inv_and.O word1.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1935 word1.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1936 a_111840_190# word1.byte2.dff_7.CLK a_111280_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1937 VDD word8.byte3.buf_RE0.O word8.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1938 a_157900_11064# a_158230_11904# a_158130_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1939 a_20820_306# word1.byte4.tinv5.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1940 word3.byte1.cgate0.inv1.I word3.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1941 a_162450_11114# a_161830_11904# a_162340_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1942 a_4660_10498# a_2820_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1943 word2.byte4.dff_3.O word2.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1944 a_17220_9714# word7.byte4.tinv4.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1945 a_166260_680# a_166050_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1946 a_66180_10088# a_65970_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1947 a_65350_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1948 VSS a_139800_1706# a_140460_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1949 a_108630_9598# word7.byte2.dff_7.CLK a_108520_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1950 word5.byte4.dff_4.O word5.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1951 VDD buf_in7.inv0.O buf_in7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1952 VDD a_103080_7976# a_104640_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1953 a_164100_4840# word4.byte1.tinv6.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X1954 buf_in2.inv1.O buf_in2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1955 VSS a_162660_11764# a_162620_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1956 a_35760_10500# word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1957 buf_in24.inv1.O buf_in24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1958 a_104080_6412# word5.byte2.dff_7.CLK a_104310_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1959 word3.byte4.dff_4.O word3.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1960 word4.byte1.dff_6.O word4.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1961 a_19060_4842# a_17220_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1962 VDD a_22980_11764# word8.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1963 VSS word6.byte3.tinv7.I a_67620_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1964 buf_in5.inv1.O buf_in5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1965 VDD a_48180_11764# word8.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1966 VDD word5.byte1.tinv7.I a_167700_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1967 word8.byte1.tinv7.O word8.byte1.tinv5.EN a_160500_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1968 VSS word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1969 VDD word1.byte4.tinv1.I a_6420_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1970 VDD a_119640_5492# word4.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1971 VSS a_12180_8628# a_12140_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1972 VSS word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1973 a_19060_1706# a_17220_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1974 a_104080_3276# word3.byte2.dff_7.CLK a_104310_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1975 a_158460_4842# a_158230_5632# a_157900_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1976 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1977 VDD word8.byte1.tinv2.I a_149700_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1978 a_47250_7362# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1979 a_124680_6578# buf_out10.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1980 VSS a_2820_306# a_4380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1981 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1982 a_58770_4842# a_58150_5632# a_58660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1983 a_13620_11112# buf_out29.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X1984 a_144340_6462# a_142500_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1985 VSS a_44580_6952# a_44540_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1986 VDD word3.byte1.tinv7.I a_167700_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1987 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1988 VDD a_119640_2356# word2.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1989 VDD word4.byte1.cgate0.nand0.B word4.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1990 VSS word4.byte4.buf_RE0.O word4.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1991 word7.byte4.dff_1.O word7.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1992 a_75360_7364# word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1993 a_100810_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1994 VDD word1.buf_ck1.I word1.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1995 VDD a_155460_6952# a_155420_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1996 a_158460_1706# a_158230_2496# a_157900_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1997 a_151650_7978# word6.byte1.dff_7.CLK a_151540_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1998 a_58770_1706# a_58150_2496# a_58660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1999 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2000 a_124680_3442# buf_out10.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2001 a_47250_4226# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2002 word4.byte1.tinv7.O buf_out7.inv0.I a_146100_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2003 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2004 a_58050_2776# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2005 a_144340_3326# a_142500_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2006 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2007 VSS a_44580_3816# a_44540_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2008 buf_sel6.inv0.O buf_sel6.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2009 VDD word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2010 a_46020_306# word1.byte3.tinv1.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2011 VDD word2.byte1.cgate0.nand0.B word2.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2012 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2013 VSS buf_out15.inv0.O buf_out15.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2014 a_20820_9714# word7.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2015 a_115440_2776# word2.byte2.dff_7.CLK a_114880_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2016 VDD a_155460_3816# a_155420_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2017 a_100810_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2018 a_75360_4228# word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2019 VDD word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2020 a_47580_7978# a_47350_8768# a_47020_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2021 VDD a_165100_7928# a_164100_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2022 a_146100_7976# word6.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2023 a_49620_306# buf_out22.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2024 word2.byte1.tinv7.O buf_out7.inv0.I a_146100_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2025 a_67620_6578# word5.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2026 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2027 VDD word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2028 a_15740_10498# word7.byte4.cgate0.inv1.O a_15570_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2029 word8.byte3.cgate0.inv1.I word8.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2030 word5.byte4.dff_1.O word5.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2031 VDD word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2032 a_8260_9048# a_6420_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2033 a_2820_306# word1.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2034 a_75360_306# word1.byte1.cgate0.nand0.B word1.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2035 a_126520_5912# a_124680_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2036 VSS buf_re.inv0.O buf_re.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2037 a_24420_6578# word5.byte4.tinv6.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2038 a_119040_6462# word5.byte2.dff_7.CLK a_118480_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2039 VDD word6.byte4.cgate0.nand0.A a_35760_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2040 VSS word1.buf_sel0.O word1.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2041 buf_in10.inv1.O buf_in10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2042 word3.byte4.dff_1.O word3.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2043 VDD buf_out25.inv0.O Do24_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2044 VSS word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2045 a_119040_3326# word3.byte2.dff_7.CLK a_118480_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2046 word5.byte1.dff_5.O word5.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2047 word6.byte1.tinv7.O word6.byte1.tinv2.EN a_149700_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2048 Do20_buf buf_out21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2049 buf_in1.inv1.O buf_in1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2050 a_22380_10498# a_22150_9548# a_21820_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2051 a_165330_1090# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2052 a_8580_8628# a_8370_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2053 VSS a_126840_10088# a_126800_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2054 word3.byte1.dff_5.O word3.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2055 a_28020_8932# word6.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2056 a_4940_2776# a_4150_2496# a_4770_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2057 VSS a_154300_11064# a_153300_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2058 word7.byte3.cgate0.inv1.I word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2059 a_144060_11114# a_143830_11904# a_143500_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2060 a_123030_7978# a_122410_8768# a_122920_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2061 a_104920_11114# a_103080_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2062 a_147100_1656# a_147430_2496# a_147330_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2063 VSS word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2064 a_19170_4842# word4.byte4.cgate0.inv1.O a_19060_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2065 a_11860_9598# a_10020_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2066 a_22150_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2067 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2068 VDD a_108840_680# a_108800_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2069 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2070 a_150700_140# a_151030_140# a_150930_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2071 VSS buf_in11.inv0.O buf_in11.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2072 VSS word7.byte1.cgate0.nand0.B a_95160_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2073 word3.buf_sel0.O buf_sel3.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X2074 VSS a_156900_4840# a_158460_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2075 a_22150_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2076 a_162620_6462# a_161830_6412# a_162450_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2077 a_61650_9048# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2078 VSS word3.byte3.tinv1.I a_46020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2079 VDD buf_in14.inv0.O buf_in14.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2080 a_56820_4840# word4.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2081 a_65250_12184# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2082 VDD word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2083 word1.byte4.tinv7.O buf_out30.inv0.I a_10020_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2084 a_143830_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2085 a_12180_10088# a_11970_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2086 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2087 VSS word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2088 buf_in28.inv0.O Di27 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2089 buf_out14.inv1.O buf_out14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2090 a_162620_3326# a_161830_3276# a_162450_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2091 a_13620_4840# buf_out29.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2092 a_56820_1704# word2.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2093 a_105240_5492# a_105030_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2094 a_107680_9548# a_108010_9548# a_107910_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2095 a_65860_7978# a_64020_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2096 a_65020_11064# word8.byte3.cgate0.inv1.O a_65250_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2097 a_51740_9598# a_50950_9548# a_51570_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2098 a_13620_1704# buf_out29.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2099 word1.byte3.dff_6.O word1.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2100 VSS a_58980_11764# a_58940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2101 a_108800_7362# word5.byte2.dff_7.CLK a_108630_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2102 VSS Di19 buf_in20.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2103 a_104920_9048# a_103080_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2104 VDD a_26580_6952# word5.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2105 word1.byte2.dff_3.O word1.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2106 VDD a_166260_680# word1.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2107 word2.byte2.tinv7.O word2.byte2.tinv0.EN a_103080_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2108 a_95160_2660# word2.byte2.cgate0.nand0.A word2.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2109 Do2_buf buf_out3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2110 word8.byte3.tinv7.O word8.byte3.tinv4.EN a_56820_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2111 VSS a_62580_5492# word4.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2112 a_1380_6952# a_1170_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2113 a_60420_7976# word6.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2114 a_108800_4226# word3.byte2.dff_7.CLK a_108630_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2115 a_104410_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2116 VSS a_159060_10088# a_159020_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2117 a_66180_8628# a_65970_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2118 VDD a_26580_3816# word3.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2119 a_103080_4840# word4.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2120 a_95160_5796# word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2121 a_160500_6578# word5.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2122 VSS word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2123 VSS a_64020_11112# a_65580_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2124 a_1380_3816# a_1170_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2125 VDD a_118480_9548# a_117480_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2126 a_162450_9598# a_161830_9548# a_162340_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2127 a_101600_7978# word6.byte2.dff_7.CLK a_101430_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2128 a_155250_7978# a_154630_8768# a_155140_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2129 buf_we3.inv0.O WE2 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X2130 VSS a_42420_6578# a_43980_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2131 word8.byte1.dff_1.O word8.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2132 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2133 VDD a_19380_8628# word6.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2134 VSS word3.byte1.nand.B a_78780_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2135 a_160500_3442# word3.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2136 VSS word5.byte2.tinv7.I a_128280_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2137 a_26370_1706# word2.byte4.cgate0.inv1.O a_26260_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2138 a_150700_7928# a_151030_8768# a_150930_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2139 word7.byte4.dff_2.O word7.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2140 VSS word8.byte2.nand.OUT word8.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2141 a_39820_4792# word4.byte3.cgate0.inv1.O a_40050_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2142 word1.byte3.cgate0.inv1.I word1.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2143 VSS a_42420_3442# a_43980_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2144 a_123240_11764# a_123030_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2145 VSS a_164100_1704# a_165660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2146 a_39820_1656# word2.byte3.cgate0.inv1.O a_40050_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2147 buf_in10.inv1.O buf_in10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2148 a_3820_11064# a_4150_11904# a_4050_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2149 VSS a_123240_11764# a_123200_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2150 a_101640_6952# a_101430_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2151 VDD a_22980_10088# word7.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2152 VDD buf_out7.inv0.I buf_out7.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X2153 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2154 VDD a_48180_10088# word7.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2155 VDD buf_in27.inv0.O buf_in27.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2156 a_101640_3816# a_101430_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2157 a_112440_2356# a_112230_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2158 VSS Di26 buf_in27.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2159 buf_in4.inv1.O buf_in4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2160 a_18780_9598# word7.byte4.cgate0.inv1.O a_18220_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2161 VDD a_122080_6412# a_121080_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2162 VSS a_66180_2356# a_66140_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2163 a_11250_9598# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2164 buf_in21.inv1.O buf_in21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2165 VDD a_65020_140# a_64020_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2166 a_64020_9714# word7.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2167 VSS A2 dec8.and4_3.nand1.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2168 word8.byte2.tinv7.O buf_out14.inv0.I a_110280_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2169 VDD a_122080_3276# a_121080_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2170 a_104310_5912# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2171 buf_sel3.inv1.O buf_sel3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2172 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2173 VDD word7.buf_sel0.O word7.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2174 word6.byte1.dff_1.O word6.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2175 a_4380_2776# word2.byte4.cgate0.inv1.O a_3820_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2176 VSS word2.byte4.tinv3.I a_13620_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2177 VDD buf_in19.inv0.O buf_in19.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2178 a_60420_11112# word8.byte3.tinv5.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2179 a_54220_140# word1.byte3.cgate0.inv1.O a_54450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2180 a_113880_306# word1.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2181 VDD A1 dec8.and4_7.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2182 a_122080_7928# word6.byte2.dff_7.CLK a_122310_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2183 VSS a_40980_8628# word6.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2184 VDD word4.byte2.tinv4.I a_117480_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2185 VDD word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2186 VDD word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2187 a_46020_9714# word7.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2188 a_7980_6462# word5.byte4.cgate0.inv1.O a_7420_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2189 a_105030_190# word1.byte2.dff_7.CLK a_104920_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2190 VSS buf_in14.inv0.O buf_in14.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2191 word4.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2192 word4.byte4.tinv7.O word4.byte4.tinv6.EN a_24420_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2193 word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.latch0.I0.O a_92280_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2194 a_65250_7978# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2195 VDD word2.byte2.tinv4.I a_117480_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2196 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2197 word5.byte4.inv_and.O word5.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2198 VSS word3.buf_ck1.I word3.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2199 VDD word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2200 VDD word4.byte1.cgate0.nand0.B word4.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2201 word4.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2202 a_7980_3326# word3.byte4.cgate0.inv1.O a_7420_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2203 VDD a_119640_5492# a_119600_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2204 a_43750_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2205 a_50950_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2206 word1.byte2.cgate0.nand0.A word1.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2207 word2.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2208 VDD word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2209 VDD a_118480_4792# a_117480_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2210 a_162060_6462# word5.byte1.dff_7.CLK a_161500_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2211 buf_in16.inv1.O buf_in16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2212 a_62370_6462# word5.byte3.cgate0.inv1.O a_62260_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2213 VDD word4.byte4.inv_and.O a_36120_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2214 a_147330_190# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2215 word2.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2216 VDD a_119640_2356# a_119600_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2217 VDD word2.byte1.cgate0.nand0.B word2.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2218 buf_out10.inv1.O buf_out10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2219 VDD a_118480_1656# a_117480_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2220 a_162060_3326# word3.byte1.dff_7.CLK a_161500_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2221 VDD a_26580_11764# a_26540_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2222 a_62370_3326# word3.byte3.cgate0.inv1.O a_62260_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2223 VSS word6.byte2.tinv5.I a_121080_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2224 VDD word2.byte4.inv_and.O a_36120_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2225 VDD word7.byte1.cgate0.nand0.B word7.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2226 Do0_buf buf_out1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2227 a_108520_7978# a_106680_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2228 a_144060_10498# a_143830_9548# a_143500_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2229 a_51460_11114# a_49620_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2230 a_51180_9598# word7.byte3.cgate0.inv1.O a_50620_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2231 a_104920_10498# a_103080_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2232 a_144660_2356# a_144450_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2233 buf_in26.inv1.O buf_in26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2234 VSS word1.byte3.buf_RE0.O word1.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2235 VSS a_48180_680# word1.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2236 VSS word1.byte1.buf_RE1.I word1.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2237 word4.byte2.dff_6.O word4.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2238 VSS a_105240_5492# word4.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2239 buf_sel1.inv0.I dec8.and4_0.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2240 VSS a_122080_7928# a_121080_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2241 VDD a_122080_11064# a_121080_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2242 a_148260_6952# a_148050_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2243 buf_sel4.inv1.O buf_sel4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2244 a_111510_2776# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2245 a_47350_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2246 VSS a_65020_1656# a_64020_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2247 word2.byte2.dff_6.O word2.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2248 word3.byte2.tinv7.O word3.byte2.tinv5.EN a_121080_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2249 VDD a_220_6412# a_120_6462# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2250 a_20820_11112# word8.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2251 a_146100_306# word1.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2252 a_158230_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2253 a_6420_7976# buf_out31.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2254 a_155420_9048# a_154630_8768# a_155250_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2255 a_148260_3816# a_148050_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2256 a_101040_2776# word2.byte2.dff_7.CLK a_100480_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2257 VDD a_150700_7928# a_149700_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2258 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2259 a_121080_6578# word5.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2260 a_47350_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2261 a_44540_4842# word4.byte3.cgate0.inv1.O a_44370_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2262 a_131700_7976# word6.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2263 VSS word7.byte3.nand.OUT word7.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2264 VDD a_220_3276# a_120_3326# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2265 a_161730_12184# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2266 a_158230_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2267 VSS word3.gt_re1.O word3.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2268 VDD word1.byte4.cgate0.nand0.A a_35760_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2269 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B a_132960_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2270 a_65020_9548# word7.byte3.cgate0.inv1.O a_65250_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2271 VDD word6.buf_ck1.I word6.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2272 a_113880_9714# buf_out13.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2273 a_44540_1706# word2.byte3.cgate0.inv1.O a_44370_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2274 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2275 VSS buf_in27.inv0.O buf_in27.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2276 a_10020_6578# word5.byte4.tinv2.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2277 a_93540_7976# word6.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2278 word8.byte3.dff_3.O word8.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2279 a_151030_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2280 a_161500_11064# word8.byte1.dff_7.CLK a_161730_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2281 a_17220_11112# word8.byte4.tinv4.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2282 a_51780_11764# a_51570_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2283 a_161830_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2284 a_150930_1090# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2285 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2286 a_11020_6412# a_11350_6412# a_11250_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2287 word2.byte2.tinv7.O word2.byte2.tinv7.EN a_128280_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2288 a_19380_680# a_19170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2289 word8.byte1.tinv7.O word8.byte1.tinv3.EN a_153300_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2290 VDD a_65020_9548# a_64020_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2291 a_121080_306# word1.byte2.tinv5.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2292 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2293 VSS word2.byte2.nand.OUT word2.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2294 a_78780_2660# buf_we2.inv1.O word2.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2295 word8.byte2.dff_1.O word8.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2296 VSS word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2297 a_128280_5796# word4.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2298 word7.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2299 a_11020_3276# a_11350_3276# a_11250_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2300 a_450_12184# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2301 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2302 a_36120_2660# word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2303 VSS word7.byte2.tinv1.I a_106680_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2304 a_42420_7976# word6.byte3.tinv0.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2305 a_58940_1090# word1.byte3.cgate0.inv1.O a_58770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2306 word4.byte2.nand.OUT buf_we3.inv1.O a_90120_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2307 word4.byte3.inv_and.O word4.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2308 a_126800_7978# word6.byte2.dff_7.CLK a_126630_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2309 a_142500_6578# buf_out8.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2310 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2311 VSS a_112440_2356# word2.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2312 VDD a_44580_8628# word6.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2313 a_123240_10088# a_123030_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2314 word4.byte4.dff_4.O word4.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2315 a_92280_7364# word5.byte2.cgate0.latch0.I0.ENB word5.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2316 VSS word1.byte1.tinv6.I a_164100_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2317 a_220_11064# word8.byte4.cgate0.inv1.O a_450_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2318 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2319 a_142500_3442# buf_out8.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2320 a_65020_4792# word4.byte3.cgate0.inv1.O a_65250_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2321 VDD word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2322 a_110280_4840# word4.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2323 VDD buf_sel6.inv0.O buf_sel6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2324 VSS a_116040_6952# word5.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2325 VDD buf_out15.inv0.I buf_out15.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X2326 a_92280_4228# word3.byte2.cgate0.latch0.I0.ENB word3.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2327 VDD word6.gt_re1.O word6.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2328 a_73020_6578# word5.byte3.cgate0.nand0.A word5.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2329 a_65020_1656# word2.byte3.cgate0.inv1.O a_65250_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2330 a_147330_6462# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2331 a_126840_6952# a_126630_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2332 a_110280_1704# word2.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2333 VDD word6.byte4.buf_RE0.O word6.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2334 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2335 VSS a_116040_3816# word3.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2336 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2337 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2338 a_51460_1090# a_49620_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2339 a_144340_5912# a_142500_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2340 buf_in12.inv1.O buf_in12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2341 VDD a_220_11064# a_120_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2342 word5.byte3.tinv7.O word5.byte3.tinv0.EN a_42420_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2343 VSS a_44580_5492# a_44540_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2344 VSS a_120_11114# a_780_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2345 a_147330_3326# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2346 a_61750_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2347 VDD word8.byte1.cgate0.nand0.B word8.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2348 a_126840_3816# a_126630_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2349 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2350 VSS buf_out30.inv0.O Do29_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2351 buf_in3.inv1.O buf_in3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2352 VDD word7.byte4.tinv6.I a_24420_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2353 VDD a_18220_7928# a_17220_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2354 buf_in26.inv1.O buf_in26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2355 VDD a_100380_4842# a_101040_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2356 VSS word4.byte4.tinv1.I a_6420_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2357 a_148050_6462# a_147430_6412# a_147940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2358 VDD a_151860_680# word1.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2359 a_160500_1704# word2.byte1.tinv5.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2360 a_61750_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2361 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2362 buf_in8.inv1.O buf_in8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2363 a_119640_8628# a_119430_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2364 a_51780_680# a_51570_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2365 a_33420_8932# word6.byte4.cgate0.nand0.A word6.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2366 VDD a_100380_1706# a_101040_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2367 a_148050_3326# a_147430_3276# a_147940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2368 word7.byte3.tinv7.O buf_out22.inv0.I a_49620_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2369 VSS a_144660_10088# a_144620_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2370 VSS word4.buf_ck1.I word4.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2371 buf_in32.inv1.O buf_in32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2372 VSS buf_in18.inv0.O buf_in18.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2373 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2374 word5.byte1.cgate0.nand0.A word5.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2375 CLK buf_ck.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2376 a_140850_7978# a_140230_8768# a_140740_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2377 word5.byte4.dff_3.O word5.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2378 a_119040_5912# word4.byte2.dff_7.CLK a_118480_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2379 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2380 word3.byte1.cgate0.nand0.A word3.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2381 a_49620_4840# word4.byte3.tinv2.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2382 VDD a_7420_4792# a_6420_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2383 word8.byte1.inv_and.O word8.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2384 word5.byte2.cgate0.inv1.I word5.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2385 VDD a_139800_6462# a_140460_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2386 a_18450_1090# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2387 a_11970_1706# word2.byte4.cgate0.inv1.O a_11860_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2388 word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.latch0.I0.ENB a_36120_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2389 a_43750_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2390 word1.byte1.tinv7.O word1.byte1.tinv5.EN a_160500_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2391 a_51740_190# a_50950_140# a_51570_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2392 word3.byte4.dff_3.O word3.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2393 VDD word5.byte3.tinv3.I a_53220_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2394 word2.byte4.dff_6.O word2.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2395 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2396 a_28020_9714# word7.byte4.tinv7.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2397 a_7980_190# word1.byte4.cgate0.inv1.O a_7420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2398 VDD a_7420_1656# a_6420_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2399 a_58050_12184# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2400 a_155140_12184# a_153300_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2401 a_55170_7978# word6.byte3.cgate0.inv1.O a_55060_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2402 word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.latch0.I0.O a_75720_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2403 word3.byte2.cgate0.inv1.I word3.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2404 VDD a_139800_3326# a_140460_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2405 a_165430_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2406 VDD a_26580_10088# a_26540_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2407 word6.byte3.dff_7.O word6.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2408 word1.byte2.tinv7.O word1.byte2.tinv1.EN a_106680_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2409 VSS a_148260_6952# word5.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2410 buf_out9.inv1.O buf_out9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2411 word5.byte4.cgate0.inv1.I word5.byte4.cgate0.nand0.A a_33420_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2412 VDD a_113880_306# a_115440_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2413 VDD word3.byte3.tinv3.I a_53220_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2414 VDD word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2415 a_12140_2776# a_11350_2496# a_11970_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2416 a_51460_10498# a_49620_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2417 VSS a_148260_3816# word3.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2418 VDD word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2419 VDD a_148260_11764# a_148220_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2420 VDD word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2421 a_151540_2776# a_149700_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2422 a_22150_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2423 a_122640_12184# word8.byte2.dff_7.CLK a_122080_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2424 a_15740_6462# a_14950_6412# a_15570_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2425 VSS a_51780_2356# a_51740_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2426 VDD word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2427 Do4_buf buf_out5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2428 a_33420_12068# word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2429 VSS a_54220_140# a_53220_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2430 VSS a_22980_8628# a_22940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2431 VDD a_50620_140# a_49620_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2432 VSS a_123240_6952# a_123200_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2433 a_162620_5912# a_161830_5632# a_162450_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2434 VSS buf_in2.inv0.O buf_in2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2435 VDD word7.byte3.buf_RE0.O word7.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2436 a_58050_7362# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2437 a_15740_3326# a_14950_3276# a_15570_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2438 dec8.and4_2.nand0.OUT dec8.and4_6.nand0.A a_67620_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2439 a_161730_4842# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2440 a_115440_7362# a_115210_6412# a_114880_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2441 VDD buf_out20.inv0.I buf_out20.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X2442 a_115830_11114# a_115210_11904# a_115720_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2443 VSS a_123240_3816# a_123200_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2444 VDD a_4980_680# a_4940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2445 a_146100_3442# word3.byte1.tinv1.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2446 a_58050_4226# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2447 a_122310_12184# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2448 word7.byte2.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2449 a_161730_1706# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2450 a_58380_1090# a_58150_140# a_57820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2451 a_142500_11112# word8.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2452 VSS buf_sel6.inv0.O buf_sel6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2453 a_107910_9048# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2454 a_115440_4226# a_115210_3276# a_114880_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2455 a_112120_9598# a_110280_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2456 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2457 word4.byte4.tinv7.O word4.byte4.tinv2.EN a_10020_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2458 a_156900_7976# word6.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2459 VSS word5.byte1.tinv1.I a_146100_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2460 VDD buf_sel1.inv0.O buf_sel1.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2461 word7.byte3.dff_3.O word7.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2462 a_50850_7978# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2463 a_60420_9714# word7.byte3.tinv5.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2464 a_122080_11064# word8.byte2.dff_7.CLK a_122310_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2465 a_161500_9548# word7.byte1.dff_7.CLK a_161730_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2466 word6.byte2.tinv7.O buf_out13.inv0.I a_113880_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2467 a_13620_6578# word5.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2468 a_14950_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2469 a_1380_5492# a_1170_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2470 a_3820_9548# a_4150_9548# a_4050_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2471 VSS buf_in32.inv0.O buf_in32.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2472 VSS a_47020_6412# a_46020_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2473 a_13620_3442# word3.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2474 buf_in10.inv1.O buf_in10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2475 word8.byte2.tinv7.O word8.byte2.tinv3.EN a_113880_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2476 VSS a_15780_10088# word7.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2477 VDD buf_re.inv1.O word8.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2478 a_4940_7362# word5.byte4.cgate0.inv1.O a_4770_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2479 VSS Di28 buf_in29.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2480 buf_re.inv1.O buf_re.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2481 a_62260_4842# a_60420_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2482 VSS a_42420_4840# a_43980_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2483 word6.byte4.cgate0.inv1.I word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2484 VSS a_47020_3276# a_46020_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2485 VDD a_155460_11764# word8.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2486 VDD a_161500_9548# a_160500_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2487 VSS word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2488 a_106680_7976# word6.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2489 VSS word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2490 VSS word1.byte2.buf_RE1.I word1.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2491 VDD RE buf_re.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2492 VSS a_1380_2356# word2.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2493 buf_in23.inv1.O buf_in23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2494 VSS a_17220_1704# a_18780_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2495 a_4940_4226# word3.byte4.cgate0.inv1.O a_4770_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2496 a_147100_6412# word5.byte1.dff_7.CLK a_147330_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2497 VDD Di3 buf_in4.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2498 a_550_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2499 a_62260_1706# a_60420_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2500 word8.byte2.tinv7.O buf_out9.inv0.I a_128280_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2501 CLK buf_ck.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2502 VDD a_162660_5492# word4.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2503 a_67620_8932# word6.byte3.tinv7.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2504 a_220_9548# word7.byte4.cgate0.inv1.O a_450_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2505 VSS a_139900_7928# a_139800_7978# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2506 VSS word1.byte4.tinv4.I a_17220_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2507 VSS a_159060_680# a_159020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2508 VSS word2.byte1.cgate0.nand0.B a_73020_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2509 a_147100_3276# word3.byte1.dff_7.CLK a_147330_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2510 VSS a_142500_9714# a_144060_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2511 a_62580_5492# a_62370_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2512 VSS a_4980_6952# word5.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2513 a_167700_7364# buf_out1.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2514 VDD A1 dec8.and4_3.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2515 a_6420_306# buf_out31.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2516 VSS a_50620_1656# a_49620_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2517 VSS word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2518 VDD a_162660_2356# word2.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2519 word4.byte3.cgate0.inv1.I word4.byte3.cgate0.nand0.A a_73020_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2520 a_131700_1092# word1.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2521 a_143830_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2522 VSS a_108840_8628# word6.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2523 a_141020_9048# a_140230_8768# a_140850_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2524 a_139900_7928# word6.byte1.dff_7.CLK a_140130_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2525 a_62580_2356# a_62370_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2526 a_167700_4228# buf_out1.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2527 VSS a_4980_3816# word3.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2528 VDD buf_sel7.inv0.O buf_sel7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2529 a_25650_11114# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2530 a_75720_7364# word5.byte3.cgate0.latch0.I0.ENB word5.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2531 VDD word1.buf_ck1.I word1.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2532 VSS word3.byte3.tinv4.I a_56820_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2533 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2534 a_143830_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2535 VDD a_220_9548# a_120_9598# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2536 a_129540_306# word1.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2537 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2538 a_93540_1092# word1.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2539 word7.byte4.tinv7.O word7.byte4.tinv5.EN a_20820_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2540 buf_in11.inv1.O buf_in11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2541 a_75720_4228# word3.byte3.cgate0.latch0.I0.ENB word3.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2542 VDD word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2543 a_118480_9548# a_118810_9548# a_118710_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2544 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2545 buf_in16.inv1.O buf_in16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2546 VSS a_111280_9548# a_110280_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2547 word5.byte3.tinv7.O word5.byte3.tinv7.EN a_67620_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2548 VDD word6.byte4.tinv6.I a_24420_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2549 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2550 VDD word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2551 VDD word7.byte1.tinv1.I a_146100_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2552 buf_in7.inv1.O buf_in7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2553 VDD a_124680_4840# a_126240_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2554 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2555 a_7980_5912# word4.byte4.cgate0.inv1.O a_7420_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2556 a_24420_11112# word8.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2557 VDD a_26580_8628# a_26540_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2558 a_15180_6462# word5.byte4.cgate0.inv1.O a_14620_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2559 VSS a_49620_1704# a_51180_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2560 word1.byte1.dff_2.O word1.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2561 VDD a_124680_1704# a_126240_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2562 a_113880_4840# word4.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2563 buf_in31.inv1.O buf_in31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2564 a_26370_6462# a_25750_6412# a_26260_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2565 a_112400_1090# word1.byte2.dff_7.CLK a_112230_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2566 VSS a_20820_7976# a_22380_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2567 VDD a_114880_11064# a_113880_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2568 word1.byte4.tinv7.O word1.byte4.tinv3.EN a_13620_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2569 VDD buf_in22.inv0.O buf_in22.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2570 a_15180_3326# word3.byte4.cgate0.inv1.O a_14620_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2571 a_162060_5912# word4.byte1.dff_7.CLK a_161500_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2572 a_166050_7978# a_165430_8768# a_165940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2573 word4.byte1.dff_0.O word4.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2574 a_62370_4842# word4.byte3.cgate0.inv1.O a_62260_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2575 word6.byte4.tinv7.O word6.byte4.tinv7.EN a_28020_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2576 VSS a_53220_6578# a_54780_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2577 a_62540_12184# a_61750_11904# a_62370_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2578 a_26370_3326# a_25750_3276# a_26260_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2579 buf_sel2.inv0.O buf_sel2.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2580 a_100810_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2581 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2582 VDD a_164100_6578# a_165660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2583 a_161500_7928# a_161830_8768# a_161730_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2584 word2.byte2.dff_4.O word2.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2585 a_126010_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2586 a_165430_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2587 VDD a_2820_306# a_4380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2588 word2.byte1.dff_0.O word2.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2589 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2590 VDD word1.gt_re1.O word1.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2591 VSS a_53220_3442# a_54780_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2592 a_50620_4792# word4.byte3.cgate0.inv1.O a_50850_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2593 word5.byte2.inv_and.O word5.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2594 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2595 VDD a_164100_3442# a_165660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2596 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2597 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2598 word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.latch0.I0.ENB a_36120_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2599 VDD word1.byte4.buf_RE0.O word1.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2600 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2601 VDD a_148260_10088# a_148220_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2602 a_50620_1656# word2.byte3.cgate0.inv1.O a_50850_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2603 VSS word3.buf_sel0.O word3.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2604 a_8540_9598# a_7750_9548# a_8370_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2605 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2606 a_112440_6952# a_112230_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2607 word3.byte2.inv_and.O word3.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2608 VDD word4.byte2.buf_RE1.I word4.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2609 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2610 VDD a_66180_6952# a_66140_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2611 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2612 buf_out13.inv1.O buf_out13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2613 word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.latch0.I0.ENB a_36120_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2614 word4.byte3.tinv7.O buf_out20.inv0.I a_56820_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2615 a_8260_12184# a_6420_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2616 VDD word2.byte2.buf_RE1.I word2.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2617 a_112440_3816# a_112230_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2618 a_148260_5492# a_148050_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2619 a_104080_140# a_104410_140# a_104310_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2620 Do3_buf buf_out4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2621 VDD a_66180_3816# a_66140_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2622 a_47350_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2623 a_4380_7362# a_4150_6412# a_3820_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2624 word2.byte3.tinv7.O buf_out20.inv0.I a_56820_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2625 VDD a_57820_9548# a_56820_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2626 VSS word2.byte1.cgate0.nand0.B a_134580_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2627 a_62370_11114# a_61750_11904# a_62260_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2628 a_22050_9598# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2629 VSS a_116040_8628# a_116000_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2630 a_115830_9598# a_115210_9548# a_115720_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2631 a_147940_9048# a_146100_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2632 buf_in29.inv1.O buf_in29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2633 word1.byte1.dff_4.O word1.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2634 word2.byte1.tinv7.O word2.byte1.tinv1.EN a_146100_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2635 VDD word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2636 a_1340_190# a_550_140# a_1170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2637 a_4380_4226# a_4150_3276# a_3820_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2638 VSS buf_out19.inv0.I buf_out19.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X2639 a_103080_11112# word8.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2640 a_1060_9598# a_120_9598# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2641 a_147430_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2642 VSS word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2643 VSS a_165100_4792# a_164100_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2644 a_146100_4840# word4.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2645 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2646 a_124680_9714# word7.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2647 word6.byte3.tinv7.O word6.byte3.tinv5.EN a_60420_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2648 VDD word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2649 dec8.and4_3.nand1.A A2 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2650 a_122080_9548# word7.byte2.dff_7.CLK a_122310_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2651 a_144620_7978# word6.byte1.dff_7.CLK a_144450_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2652 word5.byte1.tinv7.O buf_out3.inv0.I a_160500_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2653 VSS buf_sel3.inv0.O buf_sel3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2654 VSS word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2655 VSS word4.byte4.cgate0.nand0.A a_35760_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2656 word7.byte3.cgate0.nand0.A word7.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2657 buf_sel3.inv0.O buf_sel3.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2658 VSS word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2659 VSS word8.byte1.cgate0.nand0.B a_95160_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2660 a_140460_9048# word6.byte1.dff_7.CLK a_139900_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2661 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2662 VSS CLK word3.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2663 word8.byte4.dff_2.O word8.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2664 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2665 a_40770_7978# word6.byte3.cgate0.inv1.O a_40660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2666 word3.byte1.tinv7.O buf_out3.inv0.I a_160500_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2667 a_11020_4792# a_11350_5632# a_11250_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2668 a_128280_6578# word5.byte2.tinv7.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2669 VDD word8.byte3.dff_0.O_bar a_42420_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2670 word6.byte3.dff_3.O word6.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2671 buf_in16.inv1.O buf_in16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2672 a_57820_1656# a_58150_2496# a_58050_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2673 VDD word6.buf_sel0.O word6.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2674 VDD a_155460_10088# word7.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2675 a_119320_1090# a_117480_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2676 a_144660_6952# a_144450_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2677 a_1170_11114# word8.byte4.cgate0.inv1.O a_1060_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2678 a_19340_12184# a_18550_11904# a_19170_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2679 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2680 a_61980_9598# word7.byte3.cgate0.inv1.O a_61420_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2681 a_144660_3816# a_144450_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2682 a_155460_2356# a_155250_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2683 buf_in3.inv1.O buf_in3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2684 a_54550_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2685 a_111510_7362# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2686 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2687 VSS a_116040_5492# word4.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2688 VSS buf_out3.inv0.O Do2_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2689 VSS word7.byte4.dff_0.O_bar a_2820_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2690 word7.byte3.tinv7.O buf_out17.inv0.I a_67620_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2691 VDD a_24420_7976# a_25980_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2692 a_25750_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2693 VSS word6.byte1.nand.B a_39180_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2694 a_126010_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2695 VDD a_8580_11764# word8.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2696 a_101040_7362# a_100810_6412# a_100480_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2697 a_111510_4226# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2698 a_147330_5912# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2699 VDD Di31 buf_in32.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2700 buf_in18.inv0.O Di17 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2701 a_25650_10498# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2702 a_56820_1704# word2.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2703 VSS word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2704 a_43980_1090# a_43750_140# a_43420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2705 a_165100_7928# word6.byte1.dff_7.CLK a_165330_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2706 a_156900_306# word1.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2707 a_126010_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2708 a_123200_4842# word4.byte2.dff_7.CLK a_123030_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2709 a_7750_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2710 a_13620_1704# word2.byte4.tinv3.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2711 a_101040_4226# a_100810_3276# a_100480_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2712 word1.byte2.tinv7.O buf_out13.inv0.I a_113880_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2713 VSS word5.byte1.inv_and.O a_131700_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2714 a_73020_12068# word8.byte3.cgate0.nand0.A word8.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2715 a_116040_10088# a_115830_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2716 a_147940_12184# a_146100_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2717 a_147330_11114# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2718 word7.byte1.nand.B word7.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2719 a_19170_11114# a_18550_11904# a_19060_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2720 a_123200_1706# word2.byte2.dff_7.CLK a_123030_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2721 a_117480_4840# buf_out12.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2722 VDD word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2723 word7.byte3.tinv7.O word7.byte3.tinv1.EN a_46020_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2724 word5.byte2.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B a_93540_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2725 VDD word4.buf_ck1.I word4.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2726 a_161830_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2727 a_117480_1704# buf_out12.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2728 a_12180_11764# a_11970_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2729 VDD word6.byte3.tinv2.I a_49620_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2730 a_39180_6578# buf_we1.inv1.O word5.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2731 VDD word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2732 word1.byte4.cgate0.inv1.I word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2733 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2734 VDD a_143500_6412# a_142500_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2735 VSS a_146100_306# a_147660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2736 VDD word2.buf_ck1.I word2.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2737 buf_in27.inv1.O buf_in27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2738 VSS a_12180_11764# a_12140_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2739 VDD a_61420_11064# a_60420_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2740 a_154530_190# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2741 VSS word6.byte1.tinv6.I a_164100_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2742 a_146100_11112# word8.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2743 VDD a_143500_3276# a_142500_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2744 VDD a_112440_6952# word5.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2745 VSS buf_in21.inv0.O buf_in21.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2746 VDD a_146100_11112# a_147660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2747 a_100810_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2748 VDD a_118480_140# a_117480_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2749 a_126010_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2750 VSS a_46020_7976# a_47580_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2751 VDD a_55380_680# word1.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2752 VSS a_141060_6952# a_141020_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2753 VDD buf_in2.inv0.O buf_in2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2754 a_144660_680# a_144450_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2755 VDD a_112440_3816# word3.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2756 word4.byte1.dff_7.O word4.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2757 VSS a_148260_5492# word4.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2758 a_2820_306# word1.byte4.tinv0.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2759 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2760 a_10020_6578# word5.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2761 dec8.and4_3.nand1.OUT dec8.and4_3.nand1.A a_69960_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2762 word8.byte4.tinv7.O buf_out26.inv0.I a_24420_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2763 VSS a_55380_680# word1.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2764 a_154530_2776# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2765 VSS a_141060_3816# a_141020_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2766 word2.byte1.dff_7.O word2.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2767 word3.byte1.tinv7.O word3.byte1.tinv6.EN a_164100_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2768 a_11020_140# a_11350_140# a_11250_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2769 VSS word3.byte2.tinv2.I a_110280_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2770 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2771 a_144060_7978# a_143830_8768# a_143500_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2772 VDD Di16 buf_in17.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2773 a_44370_7978# a_43750_8768# a_44260_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2774 a_112230_1706# word2.byte2.dff_7.CLK a_112120_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2775 a_140850_11114# word8.byte1.dff_7.CLK a_140740_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2776 a_15740_5912# a_14950_5632# a_15570_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2777 word5.byte3.cgate0.inv1.I word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2778 VDD word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2779 a_14850_4842# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2780 a_164100_6578# word5.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2781 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2782 word6.byte3.dff_4.O word6.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2783 a_119320_190# a_117480_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2784 buf_out12.inv1.O buf_out12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2785 VSS word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2786 VDD word4.gt_re0.OUT word4.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2787 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.latch0.I0.ENB a_131700_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2788 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2789 VDD word1.byte4.tinv6.I a_24420_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2790 VSS a_123240_5492# a_123200_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2791 a_115830_6462# word5.byte2.dff_7.CLK a_115720_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2792 buf_in12.inv1.O buf_in12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2793 a_62370_9598# a_61750_9548# a_62260_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2794 VDD word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2795 a_14850_1706# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2796 word3.byte3.cgate0.inv1.I word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2797 word5.byte3.tinv7.O word5.byte3.tinv3.EN a_53220_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2798 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2799 a_166260_11764# a_166050_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2800 word6.gt_re0.OUT buf_sel6.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2801 VDD word2.gt_re0.OUT word2.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2802 VSS buf_out10.inv0.O buf_out10.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2803 a_115110_9598# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2804 a_51180_190# word1.byte3.cgate0.inv1.O a_50620_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2805 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2806 a_115830_3326# word3.byte2.dff_7.CLK a_115720_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2807 VDD a_110280_4840# a_111840_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2808 VDD a_12180_680# a_12140_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2809 VSS word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2810 Do28_buf buf_out29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2811 VDD Di5 buf_in6.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2812 VSS a_26580_11764# word8.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2813 a_104640_9598# word7.byte2.dff_7.CLK a_104080_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2814 VSS a_143500_7928# a_142500_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2815 VSS word2.byte2.tinv4.I a_117480_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2816 word8.byte2.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2817 VDD a_110280_1704# a_111840_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2818 Do29_buf buf_out30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2819 a_11970_6462# a_11350_6412# a_11860_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2820 a_151650_190# a_151030_140# a_151540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2821 word2.byte1.nand.OUT buf_we4.inv1.O a_129540_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2822 a_55060_2776# a_53220_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2823 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2824 VDD buf_out21.inv0.O Do20_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2825 word5.byte4.dff_6.O word5.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2826 VSS word7.byte1.tinv2.I a_149700_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2827 a_26260_9048# a_24420_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2828 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2829 word2.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2830 word1.byte3.cgate0.inv1.I word1.byte3.cgate0.nand0.A a_73020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2831 VSS word2.byte1.cgate0.nand0.B word2.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2832 a_4050_9048# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X2833 a_11970_3326# a_11350_3276# a_11860_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2834 VSS a_118480_1656# a_117480_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2835 VSS buf_sel4.inv0.O buf_sel4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2836 a_58660_6462# a_56820_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2837 VSS a_155460_2356# word2.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2838 word2.byte2.dff_0.O word2.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2839 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2840 a_106680_9714# word7.byte2.tinv1.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2841 VSS word2.byte4.inv_and.O a_36120_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2842 word3.byte4.dff_6.O word3.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2843 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2844 a_72300_13636# dec8.and4_4.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2845 VDD a_18220_11064# a_17220_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2846 a_165660_9048# word6.byte1.dff_7.CLK a_165100_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2847 a_12140_7362# word5.byte4.cgate0.inv1.O a_11970_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2848 a_65970_7978# word6.byte3.cgate0.inv1.O a_65860_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2849 a_8260_1090# a_6420_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2850 a_54780_4842# a_54550_5632# a_54220_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2851 a_58660_3326# a_56820_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2852 a_153300_4840# word4.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2853 a_26580_8628# a_26370_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2854 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2855 VDD word8.byte1.tinv6.I a_164100_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2856 VSS a_159060_6952# word5.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2857 VSS word7.byte3.buf_RE0.O word7.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2858 VSS a_147100_9548# a_146100_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2859 a_58980_6952# a_58770_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2860 a_12140_4226# word3.byte4.cgate0.inv1.O a_11970_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2861 a_22940_2776# a_22150_2496# a_22770_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2862 a_151540_7362# a_149700_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2863 VDD word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2864 VDD a_51780_6952# a_51740_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2865 a_54780_1706# a_54550_2496# a_54220_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2866 a_153300_1704# word2.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2867 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2868 buf_in11.inv1.O buf_in11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2869 a_8580_680# a_8370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2870 VSS a_159060_3816# word3.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2871 a_66140_9048# a_65350_8768# a_65970_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2872 VSS word1.byte2.tinv4.I a_117480_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2873 a_58980_3816# a_58770_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2874 VSS a_4980_5492# word4.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2875 VSS a_118480_11064# a_117480_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2876 a_151540_4226# a_149700_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2877 a_108240_11114# a_108010_11904# a_107680_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2878 a_2820_7976# word6.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2879 VSS a_12180_6952# word5.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2880 VDD a_51780_3816# a_51740_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2881 a_42420_7976# word6.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2882 VDD a_61420_7928# a_60420_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2883 VDD a_8580_10088# word7.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2884 VSS a_101640_8628# a_101600_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2885 VSS word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2886 VSS a_12180_3816# word3.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X2887 a_108840_5492# a_108630_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2888 VSS buf_in2.inv0.O buf_in2.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2889 word7.byte1.tinv7.O buf_out2.inv0.I a_164100_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2890 a_162660_8628# a_162450_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2891 a_15460_190# a_13620_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2892 VSS a_117480_1704# a_119040_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2893 a_6420_4840# word4.byte4.tinv1.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2894 buf_in24.inv0.O Di23 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2895 VSS word6.byte3.inv_and.O a_75720_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2896 VSS a_150700_4792# a_149700_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2897 a_131700_5796# word4.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2898 buf_in31.inv1.O buf_in31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2899 VDD buf_in17.inv0.O buf_in17.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2900 a_108840_2356# a_108630_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2901 a_147330_10498# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2902 a_108520_12184# a_106680_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2903 a_19170_9598# a_18550_9548# a_19060_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2904 VSS word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2905 VSS word4.buf_ck1.I word4.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2906 Do16_buf buf_out17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2907 a_118810_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2908 word5.byte1.cgate0.inv1.I word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2909 a_61650_1090# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2910 a_122920_9598# a_121080_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2911 VDD a_66180_5492# word4.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2912 a_93540_5796# word4.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2913 VDD buf_sel2.inv0.O buf_sel2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2914 word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.latch0.I0.O a_75720_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2915 VDD word5.gt_re1.O word5.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2916 a_12180_10088# a_11970_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X2917 a_113880_6578# word5.byte2.tinv3.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X2918 word3.byte1.cgate0.inv1.I word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2919 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2920 VDD word1.buf_sel0.O word1.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2921 VDD a_66180_2356# word2.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2922 buf_sel6.inv1.O buf_sel6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2923 a_61980_12184# word8.byte3.cgate0.inv1.O a_61420_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2924 a_15180_5912# word4.byte4.cgate0.inv1.O a_14620_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2925 a_151030_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2926 a_43420_1656# a_43750_2496# a_43650_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2927 VDD word3.gt_re1.O word3.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2928 a_53220_6578# buf_out21.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2929 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2930 VSS a_8580_2356# a_8540_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2931 VSS a_57820_6412# a_56820_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2932 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2933 VSS word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2934 VDD a_1380_6952# word5.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2935 VDD a_17220_6578# a_18780_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2936 a_75720_6578# word5.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2937 a_104920_1090# a_103080_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X2938 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2939 a_14620_7928# a_14950_8768# a_14850_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2940 a_114880_6412# a_115210_6412# a_115110_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2941 word1.byte2.tinv7.O word1.byte2.tinv3.EN a_113880_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2942 a_43420_11064# a_43750_11904# a_43650_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2943 word7.byte1.cgate0.inv1.I word7.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2944 VDD a_7420_140# a_6420_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X2945 a_53220_3442# buf_out21.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2946 VSS a_53220_4840# a_54780_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2947 VDD a_100380_11114# a_101040_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2948 VSS word5.byte1.cgate0.nand0.B a_33420_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2949 VDD a_146100_9714# a_147660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2950 VSS a_57820_3276# a_56820_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2951 VDD a_17220_3442# a_18780_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2952 VDD a_1380_3816# word3.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X2953 a_15570_9598# word7.byte4.cgate0.inv1.O a_15460_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2954 a_114880_3276# a_115210_3276# a_115110_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X2955 buf_we1.inv0.O WE0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X2956 VDD buf_in10.inv0.O buf_in10.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2957 word7.byte4.dff_7.O word7.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2958 VSS buf_in8.inv0.O buf_in8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2959 VSS buf_out21.inv0.I buf_out21.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X2960 VSS buf_in1.inv0.O buf_in1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2961 VDD a_10020_7976# a_11580_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2962 VSS a_153300_9714# a_154860_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2963 a_111610_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2964 VSS a_166260_6952# a_166220_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2965 VSS word1.buf_ck1.I word1.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2966 a_110280_1704# word2.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2967 a_1170_1706# word2.byte4.cgate0.inv1.O a_1060_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2968 VSS word8.byte4.tinv5.I a_20820_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2969 VSS word8.byte3.tinv1.I a_46020_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2970 VSS a_61420_140# a_60420_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X2971 a_150700_140# word1.byte1.dff_7.CLK a_150930_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X2972 a_7650_7978# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2973 a_36120_8932# word6.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2974 VSS word1.byte1.cgate0.nand0.B a_95160_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2975 a_101430_11114# word8.byte2.dff_7.CLK a_101320_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2976 VSS word4.gt_re1.O word4.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2977 VDD word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X2978 VSS a_166260_3816# a_166220_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2979 a_111610_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X2980 a_162450_4842# a_161830_5632# a_162340_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2981 VSS buf_ck.inv0.O CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2982 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2983 a_142500_9714# word7.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2984 a_4770_6462# word5.byte4.cgate0.inv1.O a_4660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2985 VSS a_141060_680# a_141020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2986 VSS word4.byte4.buf_RE0.O word4.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X2987 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X2988 dec8.and4_5.nand1.B A1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2989 word8.byte2.dff_7.O word8.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X2990 a_155140_9598# a_153300_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X2991 a_162450_1706# a_161830_2496# a_162340_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X2992 a_40050_4842# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X2993 VSS a_55380_10088# a_55340_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2994 a_92280_9714# word7.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X2995 VSS word7.byte2.buf_RE1.I word7.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X2996 a_103080_4840# buf_out16.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X2997 a_6420_11112# word8.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X2998 a_126840_11764# a_126630_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X2999 a_108630_7978# word6.byte2.dff_7.CLK a_108520_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3000 a_4770_3326# word3.byte4.cgate0.inv1.O a_4660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3001 VSS a_18220_4792# a_17220_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3002 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3003 buf_in11.inv1.O buf_in11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3004 VDD word1.byte3.tinv2.I a_49620_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3005 word6.byte1.tinv7.O buf_out4.inv0.I a_156900_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3006 VDD a_108840_11764# word8.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3007 VDD word6.byte2.tinv0.I a_103080_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3008 a_40050_1706# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3009 a_103080_1704# buf_out16.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3010 VDD buf_in14.inv0.I buf_in14.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3011 word8.byte1.dff_5.O word8.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3012 word5.byte4.tinv7.O buf_out29.inv0.I a_13620_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3013 a_22380_2776# word2.byte4.cgate0.inv1.O a_21820_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3014 VDD a_49620_6578# a_51180_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3015 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3016 Do27_buf buf_out28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3017 VDD a_105240_8628# a_105200_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3018 word3.byte4.tinv7.O buf_out29.inv0.I a_13620_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3019 VDD a_49620_3442# a_51180_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3020 VDD a_104080_7928# a_103080_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3021 a_25980_6462# word5.byte4.cgate0.inv1.O a_25420_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3022 a_149700_7976# word6.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3023 VSS a_7420_1656# a_6420_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3024 a_126010_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3025 VSS buf_out26.inv0.I buf_out26.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X3026 word5.byte2.dff_4.O word5.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3027 VSS word6.byte2.buf_RE1.I word6.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3028 word6.byte2.tinv7.O word6.byte2.tinv1.EN a_106680_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3029 VDD a_40980_680# word1.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3030 a_18780_12184# word8.byte4.cgate0.inv1.O a_18220_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3031 a_25980_3326# word3.byte4.cgate0.inv1.O a_25420_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3032 a_22940_11114# word8.byte4.cgate0.inv1.O a_22770_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3033 word4.byte1.dff_3.O word4.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3034 a_48140_11114# word8.byte3.cgate0.inv1.O a_47970_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3035 a_132960_9714# word7.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3036 word3.byte2.dff_4.O word3.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3037 word2.byte2.dff_7.O word2.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3038 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3039 VSS a_166260_680# a_166220_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3040 VSS word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3041 VSS word1.byte4.tinv6.I a_24420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3042 word2.byte1.dff_3.O word2.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3043 VDD EN dec8.and4_6.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3044 VSS word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3045 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3046 a_11250_12184# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3047 VSS word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3048 VSS a_65020_11064# a_64020_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3049 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.latch0.I0.ENB a_131700_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3050 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3051 word6.byte3.dff_0.O word6.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3052 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3053 a_47350_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3054 a_108240_10498# a_108010_9548# a_107680_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3055 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3056 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3057 word1.gt_re0.OUT buf_sel1.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3058 a_56820_3442# word3.byte3.tinv4.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3059 VSS word7.byte4.tinv2.I a_10020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3060 a_18220_7928# word6.byte4.cgate0.inv1.O a_18450_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3061 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3062 a_11020_11064# word8.byte4.cgate0.inv1.O a_11250_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3063 VSS word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3064 a_126010_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3065 a_119600_6462# a_118810_6412# a_119430_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3066 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3067 VSS a_6420_1704# a_7980_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3068 VSS buf_in10.inv0.O buf_in10.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3069 a_100710_9598# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3070 word7.byte2.tinv7.O buf_out10.inv0.I a_124680_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3071 a_67620_7976# word6.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3072 a_44370_190# word1.byte3.cgate0.inv1.O a_44260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3073 VSS a_126840_8628# a_126800_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3074 a_115720_4842# a_113880_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3075 buf_in6.inv1.O buf_in6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3076 a_55060_12184# a_53220_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3077 VSS word8.byte1.buf_RE1.I word8.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3078 a_119600_3326# a_118810_3276# a_119430_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3079 buf_in27.inv1.O buf_in27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3080 a_24420_7976# buf_out26.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3081 VDD word8.byte1.nand.B word8.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3082 buf_in30.inv1.O buf_in30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3083 a_40660_2776# a_39720_1706# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3084 a_118810_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3085 a_14950_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3086 a_115720_1706# a_113880_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3087 a_156900_4840# word4.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3088 VSS a_10020_11112# a_11580_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3089 a_7420_4792# word4.byte4.cgate0.inv1.O a_7650_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3090 VDD buf_in21.inv0.O buf_in21.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3091 a_36120_12068# word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3092 a_155420_1090# word1.byte1.dff_7.CLK a_155250_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3093 a_11860_9048# a_10020_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3094 VSS word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3095 word1.byte1.dff_4.O word1.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3096 word4.byte2.tinv7.O word4.byte2.tinv3.EN a_113880_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3097 a_64020_9714# buf_out18.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3098 word8.byte4.tinv7.O buf_out28.inv0.I a_17220_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3099 buf_sel4.inv0.O buf_sel4.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3100 VSS word6.byte4.tinv4.I a_17220_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3101 VSS a_141060_2356# word2.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3102 word1.byte4.tinv7.O word1.byte4.tinv5.EN a_20820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3103 VSS word1.byte3.tinv2.I a_49620_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3104 a_40980_2356# a_40770_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3105 a_7420_1656# word2.byte4.cgate0.inv1.O a_7650_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3106 VDD Di18 buf_in19.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3107 a_57820_6412# word5.byte3.cgate0.inv1.O a_58050_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3108 a_117480_6578# word5.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3109 a_450_9598# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3110 a_158850_11114# word8.byte1.dff_7.CLK a_158740_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3111 VDD word5.byte1.nand.B word5.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3112 buf_sel7.inv1.O buf_sel7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3113 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3114 a_12180_8628# a_11970_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3115 VDD word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3116 buf_out14.inv1.O buf_out14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3117 a_117480_3442# word3.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3118 a_57820_3276# word3.byte3.cgate0.inv1.O a_58050_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3119 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3120 a_33420_5796# word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3121 VDD a_100380_9598# a_101040_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3122 a_107680_7928# a_108010_8768# a_107910_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3123 a_95160_12068# word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3124 VDD word3.byte1.nand.B word3.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3125 a_155460_6952# a_155250_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3126 word4.buf_sel0.O buf_sel4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3127 word8.byte3.dff_4.O word8.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3128 a_90120_3442# word3.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3129 VDD a_146100_4840# a_147660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3130 a_54550_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3131 a_42420_306# word1.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3132 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3133 VSS a_141060_5492# a_141020_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3134 a_75720_11112# word8.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3135 a_51740_9048# a_50950_8768# a_51570_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3136 word3.byte4.tinv7.O word3.byte4.tinv4.EN a_17220_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3137 a_165100_11064# a_165430_11904# a_165330_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3138 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3139 VSS buf_in16.inv0.O buf_in16.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3140 VSS a_101640_10088# word7.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3141 VDD word4.byte3.tinv1.I a_46020_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3142 a_155460_3816# a_155250_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3143 word2.buf_sel0.O buf_sel2.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3144 VDD a_146100_1704# a_147660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3145 a_17220_6578# word5.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3146 a_54550_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3147 a_104410_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3148 VSS a_159060_8628# a_159020_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3149 a_111280_140# a_111610_140# a_111510_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3150 VDD word2.byte3.tinv1.I a_46020_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3151 word6.byte1.inv_and.O word6.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3152 VSS buf_in24.inv0.O buf_in24.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3153 VSS a_103080_1704# a_104640_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3154 VDD a_48180_5492# a_48140_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3155 VDD buf_in5.inv0.O buf_in5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3156 VSS word8.byte1.tinv0.I a_142500_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3157 word7.byte2.dff_7.O word7.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3158 VDD buf_in26.inv0.O buf_in26.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3159 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3160 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3161 VDD a_48180_2356# a_48140_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3162 a_115830_4842# word4.byte2.dff_7.CLK a_115720_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3163 buf_in22.inv1.O buf_in22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3164 VDD a_51780_5492# word4.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3165 a_167700_9714# word7.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3166 word1.byte3.tinv7.O word1.byte3.tinv1.EN a_46020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3167 VSS word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3168 word6.byte4.dff_2.O word6.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3169 VDD a_55380_11764# word8.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3170 a_6420_3442# word3.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3171 VDD a_108840_10088# word7.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3172 word7.byte2.tinv7.O word7.byte2.tinv6.EN a_124680_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3173 VSS word4.byte4.tinv6.I a_24420_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3174 a_20820_11112# buf_out27.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3175 VDD word5.byte3.buf_RE0.O word5.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3176 VDD buf_re.inv1.O word5.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3177 VDD a_51780_2356# word2.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3178 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3179 word4.byte3.nand.OUT word4.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3180 buf_sel5.inv1.O buf_sel5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3181 VDD word6.byte2.tinv7.I a_128280_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3182 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3183 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3184 VDD buf_re.inv1.O word3.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3185 VDD word3.byte3.buf_RE0.O word3.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3186 a_47580_2776# word2.byte3.cgate0.inv1.O a_47020_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3187 a_100480_6412# a_100810_6412# a_100710_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3188 word2.byte3.nand.OUT word2.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3189 VSS buf_out13.inv0.O buf_out13.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3190 word3.byte3.tinv7.O word3.byte3.tinv2.EN a_49620_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3191 a_18780_9048# word6.byte4.cgate0.inv1.O a_18220_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3192 a_11250_9048# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3193 a_58660_5912# a_56820_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3194 VDD a_25420_4792# a_24420_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3195 a_100480_3276# a_100810_3276# a_100710_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3196 a_22940_10498# word7.byte4.cgate0.inv1.O a_22770_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3197 VDD word8.buf_ck1.I word8.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3198 a_48140_10498# word7.byte3.cgate0.inv1.O a_47970_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3199 a_43650_6462# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3200 VSS buf_in29.inv0.O buf_in29.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3201 a_154530_7362# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3202 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3203 VDD a_25420_1656# a_24420_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3204 VSS a_151860_6952# a_151820_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3205 VSS a_19380_680# a_19340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3206 VSS a_159060_5492# word4.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3207 a_43650_3326# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3208 VDD buf_out24.inv0.O Do23_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3209 a_144620_11114# word8.byte1.dff_7.CLK a_144450_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3210 a_15460_7978# a_13620_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3211 a_112230_6462# a_111610_6412# a_112120_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3212 VSS word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3213 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3214 a_58980_5492# a_58770_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3215 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3216 a_2820_9714# word7.byte4.tinv0.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3217 a_154530_4226# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3218 VSS a_151860_3816# a_151820_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3219 a_55170_190# a_54550_140# a_55060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3220 VSS word2.byte2.buf_RE1.I word2.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3221 a_220_6412# a_550_6412# a_450_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3222 a_112230_3326# a_111610_3276# a_112120_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3223 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3224 a_154860_7978# a_154630_8768# a_154300_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3225 a_123030_1706# word2.byte2.dff_7.CLK a_122920_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3226 a_166220_4842# word4.byte1.dff_7.CLK a_166050_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3227 word1.byte3.dff_7.O word1.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3228 VSS a_12180_5492# word4.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3229 a_140740_9598# a_139800_9598# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3230 word2.byte3.tinv7.O word2.byte3.tinv4.EN a_56820_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3231 VSS a_40980_10088# a_40940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3232 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3233 a_15780_8628# a_15570_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3234 VSS a_161500_11064# a_160500_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3235 word1.byte1.tinv7.O buf_out4.inv0.I a_156900_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3236 a_151260_11114# a_151030_11904# a_150700_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3237 a_11020_9548# word7.byte4.cgate0.inv1.O a_11250_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3238 a_159060_10088# a_158850_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3239 VDD word1.byte2.tinv0.I a_103080_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3240 a_220_3276# a_550_3276# a_450_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3241 a_143830_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3242 a_58150_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3243 a_166220_1706# word2.byte1.dff_7.CLK a_166050_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3244 a_58150_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3245 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3246 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3247 a_131700_6578# word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3248 a_4660_4842# a_2820_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3249 buf_sel6.inv1.O buf_sel6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3250 buf_in14.inv1.O buf_in14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3251 a_55340_7978# word6.byte3.cgate0.inv1.O a_55170_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3252 word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.latch0.I0.ENB a_92280_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3253 a_101320_190# a_100380_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3254 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3255 VSS buf_in9.inv0.O buf_in9.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3256 a_125910_9598# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3257 word5.byte2.cgate0.nand0.A word5.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3258 a_4660_1706# a_2820_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3259 VDD a_117480_11112# a_119040_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3260 word6.byte4.inv_and.O word6.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3261 a_55060_7362# a_53220_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3262 VDD a_22980_680# a_22940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3263 VDD word4.buf_ck1.I word4.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3264 a_51180_9048# word6.byte3.cgate0.inv1.O a_50620_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3265 VDD a_11020_9548# a_10020_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3266 VDD buf_in12.inv0.O buf_in12.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3267 a_4980_5492# a_4770_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3268 a_108010_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3269 VSS a_153300_306# a_154860_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3270 VDD word2.buf_ck1.I word2.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3271 a_55060_4226# a_53220_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3272 buf_in26.inv0.O Di25 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3273 VSS buf_in3.inv0.O buf_in3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3274 a_65860_2776# a_64020_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3275 word5.byte2.dff_0.O word5.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3276 VDD a_155460_6952# word5.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3277 a_161730_190# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3278 a_4980_2356# a_4770_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3279 buf_in8.inv0.O Di7 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3280 a_132960_12068# word8.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3281 VDD buf_in20.inv0.O buf_in20.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3282 a_107910_1090# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3283 a_21820_9548# a_22150_9548# a_22050_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3284 a_119430_11114# word8.byte2.dff_7.CLK a_119320_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3285 VDD a_155460_3816# word3.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3286 word3.byte2.dff_0.O word3.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3287 VDD word8.byte1.buf_RE1.I word8.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3288 VSS Di17 buf_in18.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3289 a_107910_190# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3290 a_66180_2356# a_65970_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3291 a_114880_4792# a_115210_5632# a_115110_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3292 VSS word4.buf_sel0.O word4.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3293 a_22940_7362# word5.byte4.cgate0.inv1.O a_22770_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3294 word8.byte3.tinv7.O word8.byte3.tinv6.EN a_64020_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3295 a_151860_680# a_151650_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3296 word1.gt_re3.I word1.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3297 VSS word3.byte1.tinv3.I a_153300_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3298 word7.gt_re3.I word7.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3299 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3300 VSS a_62580_680# word1.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3301 a_155250_1706# word2.byte1.dff_7.CLK a_155140_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3302 a_101600_2776# a_100810_2496# a_101430_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3303 buf_sel1.inv1.O buf_sel1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3304 VDD word8.byte4.inv_and.O a_36120_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3305 a_100480_11064# a_100810_11904# a_100710_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3306 VDD word8.byte1.cgate0.nand0.B word8.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3307 VSS word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3308 VSS a_19380_6952# a_19340_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3309 VSS a_19380_2356# word2.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3310 a_22940_4226# word3.byte4.cgate0.inv1.O a_22770_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3311 a_125680_11064# a_126010_11904# a_125910_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3312 VSS a_157900_9548# a_156900_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3313 a_110280_3442# word3.byte2.tinv2.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3314 word4.byte2.tinv7.O buf_out11.inv0.I a_121080_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3315 VDD a_125680_9548# a_124680_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3316 VSS word7.byte1.cgate0.nand0.B word7.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3317 word8.byte1.dff_3.O word8.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3318 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3319 a_67620_1092# word1.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3320 a_111610_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3321 VSS a_19380_3816# a_19340_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3322 VSS a_166260_5492# a_166220_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3323 a_121080_7976# word6.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3324 a_126520_190# a_124680_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3325 a_158850_6462# word5.byte1.dff_7.CLK a_158740_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3326 VSS a_22980_6952# word5.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3327 word2.byte2.tinv7.O buf_out11.inv0.I a_121080_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3328 VSS a_126840_10088# word7.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3329 VDD word4.gt_re1.O word4.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3330 VSS word5.byte3.dff_0.O_bar a_42420_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3331 VDD a_117480_6578# a_119040_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3332 a_24420_306# buf_out26.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3333 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.latch0.I0.O a_132960_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3334 a_158130_9598# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3335 VSS word8.byte2.tinv0.I a_103080_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3336 a_158850_3326# word3.byte1.dff_7.CLK a_158740_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3337 a_10020_7976# buf_out30.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3338 VDD a_139900_140# a_139800_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3339 VSS a_22980_3816# word3.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3340 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3341 VDD word2.gt_re1.O word2.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3342 a_4770_4842# word4.byte4.cgate0.inv1.O a_4660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3343 word7.byte4.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3344 a_131700_10500# word7.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3345 VDD a_117480_3442# a_119040_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3346 VDD buf_out5.inv0.I buf_out5.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3347 VDD a_55380_10088# word7.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3348 VDD buf_in25.inv0.O buf_in25.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3349 VDD a_108840_680# word1.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3350 a_141020_1090# word1.byte1.dff_7.CLK a_140850_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3351 VDD a_54220_6412# a_53220_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3352 a_117480_1704# word2.byte2.tinv4.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3353 VSS a_149700_6578# a_151260_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3354 buf_in2.inv1.O buf_in2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3355 VSS dec8.and4_2.nand0.OUT buf_sel3.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3356 VDD word8.byte2.tinv4.I a_117480_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3357 VSS word2.buf_ck1.I word2.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3358 buf_in19.inv1.O buf_in19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3359 a_43420_6412# word5.byte3.cgate0.inv1.O a_43650_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3360 word2.byte1.dff_1.O word2.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3361 VDD a_54220_3276# a_53220_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3362 VSS a_149700_3442# a_151260_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3363 VDD a_8580_6952# a_8540_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3364 VSS word4.byte3.tinv2.I a_49620_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3365 VSS word1.buf_ck1.I word1.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3366 VSS a_57820_11064# a_56820_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3367 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3368 a_47580_11114# a_47350_11904# a_47020_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3369 a_142500_11112# buf_out8.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3370 a_122080_1656# a_122410_2496# a_122310_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3371 a_43420_140# a_43750_140# a_43650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3372 a_43420_3276# word3.byte3.cgate0.inv1.O a_43650_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3373 a_25980_5912# word4.byte4.cgate0.inv1.O a_25420_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3374 VSS a_39720_9598# a_40380_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3375 a_64020_6578# buf_out18.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3376 VDD a_8580_3816# a_8540_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3377 buf_sel2.inv1.O buf_sel2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3378 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3379 VDD word8.byte4.dff_0.O_bar a_2820_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3380 a_144620_190# a_143830_140# a_144450_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3381 a_65250_2776# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3382 VSS word3.byte3.cgate0.nand0.A a_75360_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3383 a_64020_3442# buf_out18.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3384 VDD a_1380_8628# a_1340_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3385 VDD word6.byte3.cgate0.nand0.A word6.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3386 a_47860_12184# a_46020_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3387 word7.byte2.dff_1.O word7.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3388 a_1170_6462# a_550_6412# a_1060_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3389 a_105200_11114# word8.byte2.dff_7.CLK a_105030_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3390 a_144620_10498# word7.byte1.dff_7.CLK a_144450_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3391 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3392 a_50950_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3393 VDD word8.gt_re0.OUT word8.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3394 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3395 VDD a_20820_306# a_22380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3396 VSS word1.byte2.tinv6.I a_124680_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3397 VSS a_144660_8628# a_144620_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3398 word6.byte4.tinv7.O word6.byte4.tinv0.EN a_2820_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3399 VSS buf_out29.inv0.O Do28_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3400 word6.byte3.tinv7.O buf_out24.inv0.I a_42420_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3401 a_126240_6462# word5.byte2.dff_7.CLK a_125680_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3402 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3403 a_1170_3326# a_550_3276# a_1060_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3404 VDD buf_in23.inv0.O buf_in23.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3405 VDD buf_re.inv0.O buf_re.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3406 a_108520_2776# a_106680_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3407 VDD buf_out4.inv0.O Do3_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3408 a_161500_140# word1.byte1.dff_7.CLK a_161730_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3409 a_26540_9598# a_25750_9548# a_26370_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3410 VSS word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3411 a_22660_190# a_20820_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3412 a_126240_3326# word3.byte2.dff_7.CLK a_125680_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3413 a_151260_10498# a_151030_9548# a_150700_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3414 VSS word6.byte1.cgate0.nand0.B word6.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3415 VSS word2.gt_re0.OUT word2.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3416 a_104410_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3417 VSS a_147100_140# a_146100_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3418 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.latch0.I0.O a_131700_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3419 a_119600_5912# a_118810_5632# a_119430_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3420 a_118710_4842# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3421 a_165940_9598# a_164100_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3422 VSS a_54220_7928# a_53220_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3423 word7.byte2.tinv7.O word7.byte2.tinv2.EN a_110280_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3424 word4.gt_re0.OUT buf_sel4.inv1.O a_82020_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3425 word7.byte3.cgate0.nand0.A word7.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3426 a_22380_7362# a_22150_6412# a_21820_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3427 VDD word5.byte1.cgate0.nand0.A word5.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3428 VDD word1.byte2.tinv7.I a_128280_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3429 buf_sel5.inv0.I dec8.and4_4.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3430 VDD a_39720_11114# a_40380_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3431 a_118710_1706# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3432 a_156900_6578# word5.byte1.tinv4.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3433 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3434 VDD a_117480_9714# a_119040_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3435 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3436 VDD word3.byte1.cgate0.nand0.A word3.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3437 a_22380_4226# a_22150_3276# a_21820_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3438 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3439 a_53220_11112# word8.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3440 VDD a_116040_680# a_116000_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3441 a_147940_1090# a_146100_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3442 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3443 VSS buf_in11.inv0.O buf_in11.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3444 word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.latch0.I0.ENB a_75720_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3445 a_157900_6412# a_158230_6412# a_158130_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3446 VDD a_114880_7928# a_113880_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3447 word5.byte3.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3448 a_14850_190# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3449 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3450 buf_in16.inv0.O buf_in16.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3451 a_40770_11114# word8.byte3.cgate0.inv1.O a_40660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3452 word6.byte4.cgate0.inv1.I word6.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3453 a_121080_9714# buf_out11.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3454 word1.byte2.tinv7.O word1.byte2.tinv5.EN a_121080_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3455 a_151030_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3456 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3457 a_28020_10500# word7.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3458 VSS buf_in25.inv0.O buf_in25.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3459 a_157900_3276# a_158230_3276# a_158130_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3460 buf_in7.inv0.O Di6 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3461 word5.byte2.dff_7.O word5.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3462 VDD buf_in28.inv0.O buf_in28.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3463 a_24420_11112# word8.byte4.tinv6.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3464 a_11350_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3465 a_47020_9548# a_47350_9548# a_47250_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3466 a_154630_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3467 a_47860_190# a_46020_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3468 a_153300_1704# word2.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3469 word3.byte2.dff_7.O word3.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3470 VSS buf_in31.inv0.O buf_in31.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3471 buf_in17.inv1.O buf_in17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3472 a_140460_1090# a_140230_140# a_139900_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3473 a_112120_9048# a_110280_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3474 a_40770_190# a_40150_140# a_40660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3475 a_164100_306# word1.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3476 a_11350_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3477 VSS word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3478 a_154630_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3479 a_151820_4842# word4.byte1.dff_7.CLK a_151650_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3480 word6.byte4.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3481 word1.byte3.dff_3.O word1.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3482 word6.byte2.dff_5.O word6.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3483 word8.byte2.dff_3.O word8.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3484 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3485 VSS word7.byte1.cgate0.nand0.B word7.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3486 VDD word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3487 a_126800_2776# a_126010_2496# a_126630_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3488 buf_sel2.inv1.O buf_sel2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3489 VDD a_39820_7928# a_39720_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3490 VDD a_6420_6578# a_7980_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3491 VSS a_44580_2356# word2.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3492 a_43750_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3493 word7.byte1.tinv7.O word7.byte1.tinv0.EN a_142500_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3494 a_3820_7928# a_4150_8768# a_4050_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3495 word1.byte4.cgate0.nand0.A word1.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3496 a_151820_1706# word2.byte1.dff_7.CLK a_151650_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3497 VSS word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3498 a_146100_4840# buf_out7.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3499 VSS a_61420_4792# a_60420_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3500 a_42420_4840# word4.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3501 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3502 word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.latch0.I0.ENB a_92280_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3503 VSS word7.byte4.tinv5.I a_20820_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3504 VSS a_15780_8628# word6.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3505 VDD word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3506 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3507 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3508 word1.byte4.inv_and.O word1.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3509 VDD a_6420_3442# a_7980_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3510 a_40940_7978# word6.byte3.cgate0.inv1.O a_40770_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3511 VDD word6.byte1.tinv1.I a_146100_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3512 a_146100_1704# buf_out7.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3513 VDD word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3514 VSS word5.byte3.tinv7.I a_67620_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3515 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3516 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3517 a_15460_11114# a_13620_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3518 a_40660_7362# a_39720_6462# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3519 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3520 a_40050_190# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3521 VDD buf_out13.inv0.I buf_out13.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3522 a_550_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3523 a_25750_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3524 a_146100_306# word1.byte1.tinv1.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3525 VDD a_148260_8628# a_148220_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3526 VDD word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3527 a_40660_4226# a_39720_3326# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3528 VSS buf_out4.inv0.I buf_out4.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X3529 VDD a_141060_6952# word5.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3530 word5.byte3.dff_2.O word5.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3531 VSS a_142500_7976# a_144060_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3532 a_149700_7976# word6.byte1.tinv2.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3533 a_40980_6952# a_40770_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3534 VDD buf_in6.inv0.O buf_in6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3535 VDD a_141060_3816# word3.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3536 a_119640_2356# a_119430_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3537 word3.byte3.dff_2.O word3.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3538 a_47580_10498# a_47350_9548# a_47020_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3539 a_40980_3816# a_40770_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3540 a_100480_4792# a_100810_5632# a_100710_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3541 VDD buf_out31.inv0.I buf_out31.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3542 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3543 VSS A1 dec8.and4_5.nand1.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3544 a_123240_6952# a_123030_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3545 a_140850_1706# word2.byte1.dff_7.CLK a_140740_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3546 VSS a_64020_9714# a_65580_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3547 VSS word3.byte1.buf_RE1.I word3.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3548 word7.gt_re3.I word7.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3549 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3550 a_35760_7364# word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3551 a_43650_5912# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3552 buf_sel3.inv1.O buf_sel3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3553 word8.byte4.dff_4.O word8.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3554 a_118480_7928# a_118810_8768# a_118710_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3555 a_121080_306# word1.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3556 a_123240_3816# a_123030_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3557 VSS a_151860_5492# a_151820_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3558 word5.byte1.tinv7.O word5.byte1.tinv2.EN a_149700_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3559 VSS word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3560 a_105200_10498# word7.byte2.dff_7.CLK a_105030_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3561 a_61420_7928# word6.byte3.cgate0.inv1.O a_61650_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3562 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.latch0.I0.O a_132960_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3563 a_15780_11764# a_15570_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3564 a_50950_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3565 VSS a_119640_680# a_119600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3566 a_35760_4228# word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3567 a_53220_9714# word7.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3568 VDD word4.byte3.tinv4.I a_56820_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3569 a_19340_4842# word4.byte4.cgate0.inv1.O a_19170_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3570 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3571 VDD a_103080_6578# a_104640_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3572 a_10020_306# buf_out30.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3573 a_162340_12184# a_160500_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3574 a_143730_9598# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3575 a_28020_6578# word5.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3576 VDD a_46020_306# a_47580_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3577 a_220_4792# a_550_5632# a_450_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3578 VDD word2.byte3.tinv4.I a_56820_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3579 a_19340_1706# word2.byte4.cgate0.inv1.O a_19170_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3580 VDD a_103080_3442# a_104640_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3581 a_158740_4842# a_156900_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3582 a_101430_9598# word7.byte2.dff_7.CLK a_101320_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3583 VDD word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3584 VDD a_58980_5492# a_58940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3585 word6.byte3.tinv7.O buf_out17.inv0.I a_67620_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3586 a_51570_190# word1.byte3.cgate0.inv1.O a_51460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3587 VDD buf_out26.inv0.O Do25_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3588 buf_in3.inv0.O Di2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3589 a_158740_1706# a_156900_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3590 VDD a_155460_11764# a_155420_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3591 a_103080_1704# word2.byte2.tinv0.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3592 VDD a_58980_2356# a_58940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3593 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3594 buf_in24.inv1.O buf_in24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3595 VDD a_39720_9598# a_40380_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3596 VSS word6.byte3.tinv5.I a_60420_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3597 word4.byte1.tinv7.O word4.byte1.tinv4.EN a_156900_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3598 VSS word4.byte2.tinv0.I a_103080_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3599 Do17_buf buf_out18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3600 VDD word5.byte1.tinv5.I a_160500_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3601 word1.byte1.dff_6.O word1.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3602 a_47580_7362# a_47350_6412# a_47020_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3603 dec8.and4_6.nand0.OUT dec8.and4_6.nand0.A a_74820_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3604 a_151260_4842# a_151030_5632# a_150700_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3605 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3606 a_51570_4842# a_50950_5632# a_51460_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3607 a_118480_11064# a_118810_11904# a_118710_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3608 VDD a_160500_11112# a_162060_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3609 a_17220_7976# word6.byte4.tinv4.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3610 VSS word1.byte3.tinv4.I a_56820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3611 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3612 a_8540_9048# a_7750_8768# a_8370_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3613 VDD word3.byte1.tinv5.I a_160500_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3614 a_123030_11114# a_122410_11904# a_122920_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3615 word5.byte2.tinv7.O buf_out12.inv0.I a_117480_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3616 VDD word5.byte1.nand.OUT word5.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3617 word4.byte3.dff_6.O word4.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3618 VSS word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3619 VDD a_3820_7928# a_2820_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3620 a_47580_4226# a_47350_3276# a_47020_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3621 a_44260_9598# a_42420_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3622 word1.byte2.dff_2.O word1.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3623 a_151260_1706# a_151030_2496# a_150700_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3624 VSS a_104080_4792# a_103080_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3625 a_51570_1706# a_50950_2496# a_51460_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3626 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3627 VDD word1.byte3.cgate0.nand0.A word1.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3628 a_50850_2776# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3629 word2.byte3.dff_6.O word2.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3630 VDD word3.byte1.nand.OUT word3.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3631 word3.byte2.tinv7.O buf_out12.inv0.I a_117480_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3632 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3633 a_40380_7978# a_40150_8768# a_39820_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3634 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3635 a_22050_9048# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3636 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3637 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3638 a_4150_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3639 a_122310_6462# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3640 VDD buf_in15.inv0.O buf_in15.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3641 VSS a_144660_10088# word7.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3642 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3643 VDD word4.buf_sel0.O word4.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3644 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3645 a_60420_6578# word5.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3646 word1.byte3.tinv7.O buf_out24.inv0.I a_42420_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3647 a_44580_10088# a_44370_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3648 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3649 VSS buf_in6.inv0.O buf_in6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3650 word7.byte4.tinv7.O buf_out29.inv0.I a_13620_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3651 a_149700_9714# word7.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3652 VSS buf_in27.inv0.O buf_in27.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3653 a_1060_9048# a_120_7978# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3654 a_26260_1090# a_24420_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3655 a_111840_6462# word5.byte2.dff_7.CLK a_111280_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3656 a_122310_3326# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3657 a_147430_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3658 a_4050_1090# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3659 VDD word2.buf_sel0.O word2.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3660 VDD a_8580_5492# word4.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3661 word8.byte2.tinv7.O word8.byte2.tinv5.EN a_121080_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3662 a_17220_306# word1.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3663 VSS a_19380_5492# a_19340_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3664 a_123030_6462# a_122410_6412# a_122920_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3665 a_165660_1090# a_165430_140# a_165100_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3666 a_111840_3326# word3.byte2.dff_7.CLK a_111280_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3667 VDD a_8580_2356# word2.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3668 a_65970_190# a_65350_140# a_65860_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3669 VDD a_162660_11764# word8.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3670 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3671 a_26580_680# a_26370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3672 a_123030_3326# a_122410_3276# a_122920_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3673 a_158850_4842# word4.byte1.dff_7.CLK a_158740_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3674 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3675 VDD Di1 buf_in2.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3676 VSS word8.byte4.tinv1.I a_6420_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3677 VDD EN dec8.and4_3.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3678 VSS a_22980_5492# word4.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3679 a_20820_7976# word6.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3680 word1.byte3.tinv7.O word1.byte3.tinv3.EN a_53220_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3681 word7.byte1.tinv7.O word7.byte1.tinv7.EN a_167700_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3682 a_67620_5796# word4.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3683 VSS word7.byte2.tinv3.I a_113880_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3684 a_66140_1090# word1.byte3.cgate0.inv1.O a_65970_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3685 word3.byte4.tinv7.O word3.byte4.tinv1.EN a_6420_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3686 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3687 a_15460_10498# a_13620_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3688 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3689 a_139900_1656# a_140230_2496# a_140130_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3690 VSS a_106680_9714# a_108240_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3691 a_24420_4840# word4.byte4.tinv6.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3692 VSS a_154300_6412# a_153300_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3693 VDD word7.buf_ck1.I word7.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3694 word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.latch0.I0.ENB a_75720_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3695 VDD word8.byte4.cgate0.nand0.A word8.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3696 word5.gt_re1.O word5.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3697 VDD a_101640_680# a_101600_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3698 VSS word3.byte3.buf_RE0.O word3.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3699 a_40150_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3700 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3701 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3702 VDD CLK word4.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3703 a_128280_7976# buf_out9.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3704 VDD word5.byte4.tinv7.I a_28020_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3705 a_65860_7362# a_64020_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3706 word1.byte4.cgate0.inv1.I word1.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3707 VSS a_149700_4840# a_151260_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3708 a_61980_9048# word6.byte3.cgate0.inv1.O a_61420_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3709 VSS a_154300_3276# a_153300_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3710 a_143500_6412# a_143830_6412# a_143730_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3711 VSS a_123240_6952# word5.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3712 word3.gt_re1.O word3.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3713 a_118810_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3714 VDD CLK word2.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3715 a_65860_4226# a_64020_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3716 VDD word3.byte4.tinv7.I a_28020_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3717 buf_in9.inv1.O buf_in9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3718 VSS a_43420_9548# a_42420_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3719 a_143500_3276# a_143830_3276# a_143730_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3720 VSS a_123240_3816# word3.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X3721 VSS word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3722 a_66180_6952# a_65970_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3723 VDD buf_out6.inv0.O Do5_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3724 VDD a_56820_4840# a_58380_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3725 VDD word8.byte2.inv_and.O a_92280_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3726 VDD word7.byte1.tinv3.I a_153300_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3727 buf_in5.inv1.O buf_in5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3728 a_101600_7362# word5.byte2.dff_7.CLK a_101430_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3729 VSS a_26580_2356# a_26540_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3730 a_66180_3816# a_65970_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3731 a_155250_6462# a_154630_6412# a_155140_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3732 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3733 VDD a_19380_6952# word5.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3734 VDD a_56820_1704# a_58380_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3735 VSS a_26580_680# a_26540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3736 VSS word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3737 a_116040_8628# a_115830_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3738 buf_in20.inv1.O buf_in20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3739 a_8540_11114# word8.byte4.cgate0.inv1.O a_8370_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3740 word7.byte4.dff_4.O word7.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3741 VDD a_25420_140# a_24420_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3742 VSS word6.byte1.cgate0.nand0.B a_95160_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3743 word2.buf_sel0.O buf_sel2.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X3744 a_155250_3326# a_154630_3276# a_155140_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3745 a_101600_4226# word3.byte2.dff_7.CLK a_101430_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3746 a_166050_1706# word2.byte1.dff_7.CLK a_165940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3747 VDD a_19380_3816# word3.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3748 VDD a_56820_11112# a_58380_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3749 VSS word2.byte3.tinv1.I a_46020_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3750 a_121080_3442# word3.byte2.tinv5.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3751 a_14620_140# word1.byte4.cgate0.inv1.O a_14850_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3752 VDD word1.byte1.tinv1.I a_146100_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3753 dec8.and4_5.nand0.OUT A0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3754 VSS word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3755 a_126240_5912# word4.byte2.dff_7.CLK a_125680_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3756 word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.latch0.I0.ENB a_92280_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3757 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3758 VSS buf_sel5.inv0.O buf_sel5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3759 a_46020_11112# word8.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3760 VDD word6.byte1.inv_and.O a_131700_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3761 VDD word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3762 VSS word5.byte2.tinv5.I a_121080_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3763 a_7750_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3764 a_65350_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3765 word3.gt_re3.I word3.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3766 word7.byte4.dff_0.O word7.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3767 a_25650_7978# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3768 word8.byte2.nand.OUT buf_we3.inv1.O a_90120_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3769 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3770 VDD word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3771 a_58770_11114# word8.byte3.cgate0.inv1.O a_58660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3772 word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.latch0.I0.O a_93540_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3773 word8.byte3.nand.OUT word8.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3774 VDD a_116040_11764# a_116000_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3775 VDD a_155460_10088# a_155420_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3776 a_126630_9598# word7.byte2.dff_7.CLK a_126520_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3777 a_22770_6462# word5.byte4.cgate0.inv1.O a_22660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3778 VDD buf_we1.inv1.O word6.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3779 buf_out11.inv1.O buf_out11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3780 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3781 VDD a_121080_7976# a_122640_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3782 a_22770_3326# word3.byte4.cgate0.inv1.O a_22660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3783 word5.byte1.dff_1.O word5.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3784 VSS word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3785 a_144060_190# word1.byte1.dff_7.CLK a_143500_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3786 Do1_buf buf_out2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3787 word1.byte4.dff_4.O word1.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3788 Do23_buf buf_out24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3789 a_122080_6412# word5.byte2.dff_7.CLK a_122310_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3790 VSS word2.byte1.nand.B a_78780_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3791 a_11580_9598# word7.byte4.cgate0.inv1.O a_11020_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3792 VDD a_160500_9714# a_162060_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3793 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3794 word3.byte1.dff_1.O word3.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3795 VSS word4.byte2.tinv7.I a_128280_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3796 buf_in31.inv0.O Di30 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3797 a_123030_9598# a_122410_9548# a_122920_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3798 a_108630_190# a_108010_140# a_108520_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3799 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3800 VDD a_1380_11764# a_1340_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3801 a_122080_3276# word3.byte2.dff_7.CLK a_122310_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3802 a_157900_4792# a_158230_5632# a_158130_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3803 VSS buf_out17.inv0.I buf_out17.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X3804 a_110280_11112# word8.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3805 a_65250_7362# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3806 a_162340_6462# a_160500_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3807 VSS a_62580_6952# a_62540_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3808 a_144620_2776# a_143830_2496# a_144450_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3809 buf_sel2.inv1.O buf_sel2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3810 VSS word8.byte3.inv_and.O a_75720_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3811 a_10020_7976# word6.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3812 VSS a_25420_1656# a_24420_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3813 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3814 a_153300_3442# word3.byte1.tinv3.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3815 a_65250_4226# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3816 word4.byte1.tinv7.O buf_out2.inv0.I a_164100_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3817 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3818 a_162340_3326# a_160500_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3819 a_1170_190# word1.byte4.cgate0.inv1.O a_1060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3820 VSS a_62580_3816# a_62540_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3821 VDD word4.byte2.tinv2.I a_110280_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3822 VSS buf_sel6.inv0.O buf_sel6.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3823 a_115110_9048# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3824 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3825 VSS buf_in14.inv0.O buf_in14.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3826 a_154630_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3827 a_65580_7978# a_65350_8768# a_65020_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3828 a_105240_680# a_105030_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3829 a_164100_7976# word6.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3830 VSS word7.byte4.nand.OUT word7.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3831 word2.byte1.tinv7.O buf_out2.inv0.I a_164100_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3832 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3833 a_108520_7362# a_106680_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3834 VDD word2.byte2.tinv2.I a_110280_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3835 a_104640_9048# word6.byte2.dff_7.CLK a_104080_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3836 word1.byte3.tinv7.O buf_out17.inv0.I a_67620_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3837 VDD word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3838 VSS word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3839 VDD a_112440_5492# a_112400_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3840 VDD a_111280_4792# a_110280_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3841 a_42420_6578# word5.byte3.tinv0.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3842 word6.byte3.tinv7.O buf_out21.inv0.I a_53220_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3843 VDD a_123240_11764# word8.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3844 VDD a_162660_10088# word7.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3845 a_108520_4226# a_106680_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3846 a_105200_9598# a_104410_9548# a_105030_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3847 VDD word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3848 VDD a_112440_2356# a_112400_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3849 VDD a_111280_1656# a_110280_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3850 a_26540_12184# a_25750_11904# a_26370_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3851 VDD word7.byte3.tinv2.I a_49620_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3852 VSS word1.byte4.tinv1.I a_6420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3853 buf_in20.inv1.O buf_in20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3854 VSS Di7 buf_in8.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3855 a_101320_7978# a_100380_7978# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3856 buf_we2.inv0.O WE1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X3857 buf_in1.inv1.O buf_in1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3858 VSS a_24420_1704# a_25980_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3859 a_46020_7976# word6.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3860 word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.latch0.I0.O a_92280_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3861 VDD word7.byte3.cgate0.nand0.A a_75360_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3862 VSS word7.byte1.buf_RE1.I word7.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3863 VDD a_120_7978# a_780_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3864 VSS word2.buf_ck1.I word2.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3865 word4.byte4.inv_and.O word4.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3866 word5.byte2.tinv7.O buf_out16.inv0.I a_103080_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3867 a_165100_1656# a_165430_2496# a_165330_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3868 VDD A0 dec8.and4_6.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3869 word8.byte1.nand.B word8.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3870 VDD word5.byte2.cgate0.nand0.A word5.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3871 a_141060_6952# a_140850_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3872 a_40150_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3873 word4.byte3.dff_2.O word4.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3874 VDD a_126840_680# a_126800_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3875 a_6420_11112# buf_out31.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3876 a_151030_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3877 a_50620_140# a_50950_140# a_50850_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3878 word3.byte2.tinv7.O buf_out16.inv0.I a_103080_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3879 a_141060_3816# a_140850_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3880 VDD word3.byte2.cgate0.nand0.A word3.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3881 a_25420_4792# word4.byte4.cgate0.inv1.O a_25650_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3882 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3883 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3884 a_154530_11114# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X3885 a_40150_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3886 a_26370_11114# a_25750_11904# a_26260_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3887 a_33420_306# word1.byte4.cgate0.nand0.A word1.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3888 VSS word3.byte3.tinv6.I a_64020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3889 a_33420_6578# word5.byte4.cgate0.nand0.A word5.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3890 a_151030_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3891 a_161830_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3892 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3893 a_151820_190# a_151030_140# a_151650_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3894 a_25420_1656# word2.byte4.cgate0.inv1.O a_25650_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3895 word7.byte1.dff_2.O word7.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3896 VDD word7.byte2.tinv3.I a_113880_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3897 buf_in13.inv1.O buf_in13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3898 a_11860_1090# a_10020_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3899 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3900 a_123240_5492# a_123030_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3901 VDD buf_out28.inv0.O Do27_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3902 a_125680_9548# a_126010_9548# a_125910_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X3903 a_44580_11764# a_44370_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3904 a_8540_10498# word7.byte4.cgate0.inv1.O a_8370_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3905 word1.byte4.tinv7.O word1.byte4.tinv0.EN a_2820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3906 a_75720_306# word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3907 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3908 buf_in25.inv1.O buf_in25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3909 VDD a_107680_6412# a_106680_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3910 a_126800_7362# word5.byte2.dff_7.CLK a_126630_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3911 a_122920_9048# a_121080_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3912 VDD a_44580_6952# word5.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3913 VDD a_56820_9714# a_58380_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3914 word2.byte2.tinv7.O word2.byte2.tinv5.EN a_121080_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3915 a_12180_680# a_11970_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3916 Do19_buf buf_out20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3917 a_153300_11112# word8.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3918 a_126800_4226# word3.byte2.dff_7.CLK a_126630_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3919 VDD a_107680_3276# a_106680_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3920 a_122410_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3921 a_107680_140# word1.byte2.dff_7.CLK a_107910_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X3922 VDD a_44580_3816# word3.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3923 a_121080_4840# word4.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3924 VSS buf_in19.inv0.O buf_in19.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3925 VDD a_153300_11112# a_154860_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3926 VSS word6.byte3.nand.OUT word6.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3927 word7.byte1.tinv7.O word7.byte1.tinv3.EN a_153300_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3928 VSS word2.gt_re1.O word2.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3929 VSS a_154300_140# a_153300_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3930 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B a_132960_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3931 a_119430_4842# a_118810_5632# a_119320_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3932 a_51740_1090# word1.byte3.cgate0.inv1.O a_51570_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3933 VDD a_100480_7928# a_100380_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X3934 VSS a_60420_6578# a_61980_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3935 VSS word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3936 a_10020_4840# word4.byte4.tinv2.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X3937 a_128280_1092# buf_out9.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3938 a_144060_2776# word2.byte1.dff_7.CLK a_143500_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3939 VDD word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3940 a_167700_11112# word8.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3941 VDD a_116040_10088# a_116000_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3942 a_119430_1706# a_118810_2496# a_119320_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3943 a_44370_1706# word2.byte3.cgate0.inv1.O a_44260_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3944 a_113880_7976# buf_out13.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X3945 VDD word5.byte4.tinv3.I a_13620_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3946 word2.byte3.dff_4.O word2.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3947 a_104410_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3948 VDD a_159060_680# a_159020_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3949 VSS a_60420_3442# a_61980_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3950 a_15570_7978# word6.byte4.cgate0.inv1.O a_15460_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3951 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3952 a_108240_7978# a_108010_8768# a_107680_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X3953 a_147660_6462# word5.byte1.dff_7.CLK a_147100_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3954 word6.byte4.dff_7.O word6.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3955 a_47970_6462# word5.byte3.cgate0.inv1.O a_47860_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3956 a_24420_3442# word3.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3957 VDD word3.byte4.tinv3.I a_13620_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3958 VDD word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3959 a_140130_6462# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3960 buf_out10.inv1.O buf_out10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3961 a_119640_6952# a_119430_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3962 a_75720_7976# word6.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X3963 word5.byte3.dff_5.O word5.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3964 VSS a_153300_7976# a_154860_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3965 VDD buf_in6.inv0.O buf_in6.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3966 a_22050_190# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3967 a_147660_3326# word3.byte1.dff_7.CLK a_147100_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3968 VDD word6.byte1.cgate0.nand0.B word6.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3969 a_47970_3326# word3.byte3.cgate0.inv1.O a_47860_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3970 VSS word6.byte2.tinv1.I a_106680_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3971 word1.byte4.dff_2.O word1.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3972 VDD word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3973 a_140130_3326# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3974 VDD a_1380_10088# a_1340_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3975 a_119640_3816# a_119430_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3976 word3.byte3.dff_5.O word3.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X3977 buf_in30.inv0.O Di29 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X3978 VDD a_11020_7928# a_10020_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X3979 a_140850_6462# a_140230_6412# a_140740_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3980 a_48140_6462# a_47350_6412# a_47970_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3981 VDD buf_in30.inv0.O buf_in30.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3982 Do26_buf buf_out27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X3983 a_155140_9048# a_153300_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3984 a_12180_680# a_11970_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X3985 VSS a_55380_8628# a_55340_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X3986 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X3987 a_140850_3326# a_140230_3276# a_140740_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X3988 word4.byte2.dff_2.O word4.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3989 VSS a_11020_11064# a_10020_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3990 VSS a_107680_7928# a_106680_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X3991 a_48140_3326# a_47350_3276# a_47970_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3992 a_122310_5912# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X3993 word6.byte1.dff_6.O word6.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3994 a_73020_5796# word4.byte3.cgate0.nand0.A word4.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X3995 VDD buf_out19.inv0.O Do18_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3996 VDD word1.byte1.inv_and.O a_131700_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X3997 word2.byte2.dff_2.O word2.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X3998 a_111840_5912# word4.byte2.dff_7.CLK a_111280_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X3999 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4000 a_18780_1090# a_18550_140# a_18220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4001 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4002 VDD word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4003 buf_sel8.inv0.O buf_sel8.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4004 a_11250_1090# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4005 a_117480_306# word1.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4006 a_64020_9714# word7.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4007 VSS word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4008 a_106680_6578# word5.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4009 word4.byte3.tinv7.O word4.byte3.tinv0.EN a_42420_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4010 VDD a_25420_11064# a_24420_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4011 VSS word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4012 word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.latch0.I0.O a_93540_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4013 VDD a_123240_10088# word7.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4014 a_20820_9714# word7.byte4.tinv5.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4015 VDD buf_we1.inv1.O word1.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4016 VDD word8.byte1.cgate0.nand0.B word8.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4017 VSS buf_in16.inv0.I buf_in16.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4018 a_67620_6578# word5.byte3.tinv7.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4019 VSS a_101640_680# a_101600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4020 VSS word1.gt_re1.O word1.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4021 buf_in9.inv1.O buf_in9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4022 VSS a_48180_10088# word7.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4023 VSS a_125680_11064# a_124680_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4024 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4025 a_10020_9714# buf_out30.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4026 a_115440_11114# a_115210_11904# a_114880_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4027 a_148220_12184# a_147430_11904# a_148050_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4028 a_22660_4842# a_20820_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4029 buf_in24.inv1.O buf_in24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4030 a_126520_7978# a_124680_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4031 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4032 a_162660_2356# a_162450_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4033 a_49620_11112# word8.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4034 Do25_buf buf_out26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4035 a_22660_1706# a_20820_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4036 a_143500_4792# a_143830_5632# a_143730_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4037 buf_in22.inv0.O Di21 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4038 VDD word7.byte3.buf_RE0.O word7.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4039 a_28020_8932# word6.byte4.tinv7.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4040 a_50850_7362# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4041 a_10020_306# word1.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4042 VSS a_123240_5492# word4.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4043 buf_sel2.inv0.I dec8.and4_1.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4044 word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.latch0.I0.O a_75720_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4045 a_22980_5492# a_22770_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4046 word5.byte2.tinv7.O buf_out9.inv0.I a_128280_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4047 a_166260_6952# a_166050_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4048 dec8.and4_1.nand0.OUT A0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4049 a_115720_12184# a_113880_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4050 a_115110_11114# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4051 a_154530_10498# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4052 VSS a_114880_4792# a_113880_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4053 a_26370_9598# a_25750_9548# a_26260_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4054 a_65350_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4055 a_50850_4226# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4056 word4.byte4.cgate0.inv1.I word4.byte4.cgate0.nand0.A a_33420_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4057 a_7980_11114# a_7750_11904# a_7420_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4058 VDD buf_we2.inv1.O word5.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4059 VDD word5.byte2.nand.OUT word5.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4060 a_51180_1090# a_50950_140# a_50620_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4061 a_164100_306# word1.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4062 a_22980_2356# a_22770_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4063 VSS word3.byte1.buf_RE1.I word3.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4064 word3.byte2.tinv7.O buf_out9.inv0.I a_128280_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4065 a_100710_9048# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4066 a_166260_3816# a_166050_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4067 word7.gt_re3.I word7.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4068 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4069 VDD buf_sel5.inv0.O buf_sel5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4070 VDD word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4071 a_36120_7364# word5.byte4.cgate0.latch0.I0.ENB word5.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4072 a_65350_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4073 a_62540_4842# word4.byte3.cgate0.inv1.O a_62370_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4074 a_19170_7978# a_18550_8768# a_19060_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4075 word3.byte1.nand.B word3.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4076 VDD buf_we2.inv1.O word3.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4077 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4078 VDD word3.byte2.nand.OUT word3.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4079 a_44580_10088# a_44370_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4080 word1.byte3.tinv7.O buf_out21.inv0.I a_53220_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4081 VDD a_108840_11764# a_108800_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4082 a_55380_10088# a_55170_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4083 VSS a_126840_680# a_126800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4084 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4085 a_62540_1706# word2.byte3.cgate0.inv1.O a_62370_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4086 a_36120_4228# word3.byte4.cgate0.latch0.I0.ENB word3.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4087 a_56820_4840# buf_out20.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4088 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4089 VDD a_156900_7976# a_158460_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4090 a_115210_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4091 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4092 a_144450_9598# word7.byte1.dff_7.CLK a_144340_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4093 word5.byte4.tinv7.O word5.byte4.tinv7.EN a_28020_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4094 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4095 a_141060_11764# a_140850_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4096 a_56820_1704# buf_out20.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4097 a_50620_11064# a_50950_11904# a_50850_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4098 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4099 buf_in8.inv1.O buf_in8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4100 a_115210_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4101 VSS a_141060_11764# a_141020_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4102 buf_in29.inv1.O buf_in29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4103 VDD a_153300_9714# a_154860_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4104 a_146100_1704# word2.byte1.tinv1.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4105 a_8370_4842# a_7750_5632# a_8260_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4106 word6.byte2.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4107 a_105240_8628# a_105030_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4108 a_450_9048# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4109 VDD buf_we4.inv0.O buf_we4.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4110 a_139900_6412# word5.byte1.dff_7.CLK a_140130_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4111 VSS a_10020_1704# a_11580_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4112 word2.byte2.dff_7.CLK word2.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4113 VSS word4.byte1.tinv1.I a_146100_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4114 a_8370_1706# a_7750_2496# a_8260_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4115 CLK buf_ck.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4116 a_128280_11112# word8.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4117 a_7650_2776# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4118 VSS word7.byte2.tinv6.I a_124680_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4119 a_60420_7976# word6.byte3.tinv5.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4120 a_139900_3276# word3.byte1.dff_7.CLK a_140130_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4121 a_22770_4842# word4.byte4.cgate0.inv1.O a_22660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4122 VSS word8.byte3.tinv3.I a_53220_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4123 a_160500_6578# buf_out3.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4124 VDD a_62580_8628# word6.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4125 VSS word1.byte1.buf_RE1.I word1.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4126 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4127 VSS a_101640_8628# word6.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4128 a_160500_3442# buf_out3.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4129 VSS a_24420_306# a_25980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4130 VDD a_147100_4792# a_146100_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4131 VDD word8.byte3.tinv7.I a_67620_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4132 buf_in9.inv1.O buf_in9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4133 a_49620_3442# word3.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4134 a_165330_6462# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4135 VDD word4.byte1.nand.B word4.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4136 VDD a_116040_11764# word8.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4137 VDD a_26580_6952# a_26540_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4138 VDD a_147100_1656# a_146100_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4139 a_111280_9548# a_111610_9548# a_111510_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4140 VDD buf_in12.inv0.I buf_in12.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4141 a_162340_5912# a_160500_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4142 word4.byte4.tinv7.O buf_out28.inv0.I a_17220_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4143 word5.byte3.tinv7.O word5.byte3.tinv5.EN a_60420_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4144 VSS a_62580_5492# a_62540_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4145 VSS a_105240_2356# a_105200_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4146 a_165330_3326# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4147 a_93540_11112# word8.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4148 VDD word2.byte1.nand.B word2.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4149 VSS Di2 buf_in3.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4150 VDD a_26580_3816# a_26540_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4151 Do25_buf buf_out26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4152 a_17220_7976# word6.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4153 a_166050_6462# a_165430_6412# a_165940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4154 word2.byte4.tinv7.O buf_out28.inv0.I a_17220_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4155 a_24420_306# word1.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4156 word8.byte1.cgate0.nand0.A word8.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4157 a_54450_9598# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4158 buf_in20.inv1.O buf_in20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4159 Do7_buf buf_out8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4160 VSS a_108840_6952# a_108800_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4161 a_166050_3326# a_165430_3276# a_165940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4162 VSS a_162660_10088# a_162620_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4163 VSS buf_out18.inv0.O Do17_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4164 VSS word2.byte3.tinv4.I a_56820_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4165 a_25980_12184# word8.byte4.cgate0.inv1.O a_25420_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4166 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4167 a_105030_4842# a_104410_5632# a_104920_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4168 VSS a_108840_3816# a_108800_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4169 a_55340_11114# word8.byte3.cgate0.inv1.O a_55170_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4170 word6.byte4.tinv7.O word6.byte4.tinv5.EN a_20820_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4171 VSS word7.byte1.tinv4.I a_156900_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4172 a_113880_306# buf_out13.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4173 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4174 a_6420_4840# word4.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4175 VSS buf_sel1.inv0.O buf_sel1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4176 a_104310_7978# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4177 a_105030_1706# a_104410_2496# a_104920_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4178 word7.byte4.cgate0.nand0.A word7.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4179 word4.byte3.tinv7.O word4.byte3.tinv7.EN a_67620_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4180 VDD a_147100_11064# a_146100_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4181 word2.byte3.dff_0.O word2.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4182 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4183 VDD a_144660_680# a_144620_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4184 a_46020_9714# word7.byte3.tinv1.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4185 a_6420_1704# word2.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4186 a_75720_1092# word1.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4187 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4188 VDD word7.byte2.tinv1.I a_106680_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4189 word5.byte2.dff_3.O word5.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4190 VSS a_166260_6952# word5.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4191 buf_in15.inv1.O buf_in15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4192 a_115440_10498# a_115210_9548# a_114880_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4193 a_18220_1656# a_18550_2496# a_18450_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4194 a_54550_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4195 a_1340_9598# a_550_9548# a_1170_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4196 VSS word5.byte1.nand.B a_39180_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4197 VDD word1.byte1.cgate0.nand0.B word1.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4198 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4199 a_4660_190# a_2820_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4200 VSS a_166260_3816# word3.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4201 word3.byte2.dff_3.O word3.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4202 word4.byte3.tinv7.O buf_out22.inv0.I a_49620_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4203 a_131700_10500# word7.byte1.cgate0.latch0.I0.ENB word7.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4204 a_141060_5492# a_140850_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4205 VDD word7.byte4.nand.OUT word7.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4206 a_35760_306# word1.byte1.cgate0.nand0.B word1.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4207 a_47860_4842# a_46020_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4208 a_40150_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4209 a_49620_306# word1.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4210 word2.byte3.tinv7.O buf_out22.inv0.I a_49620_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4211 buf_in4.inv1.O buf_in4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4212 word8.byte4.tinv7.O word8.byte4.tinv2.EN a_10020_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4213 a_62260_12184# a_60420_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4214 VSS a_3820_4792# a_2820_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4215 buf_in25.inv1.O buf_in25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4216 a_14950_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4217 a_144620_7362# word5.byte1.dff_7.CLK a_144450_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4218 a_115110_10498# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4219 a_140740_9048# a_139800_7978# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4220 a_47860_1706# a_46020_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4221 VSS a_40980_8628# a_40940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4222 a_159060_8628# a_158850_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4223 dec8.and4_3.nand0.OUT A0 a_69420_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4224 a_7980_10498# a_7750_9548# a_7420_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4225 VDD word7.byte4.buf_RE0.O word7.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4226 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4227 a_58150_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4228 a_48180_5492# a_47970_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4229 word1.byte3.inv_and.O word1.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4230 a_144620_4226# word3.byte1.dff_7.CLK a_144450_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4231 VSS a_42420_11112# a_43980_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4232 a_140230_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4233 VDD buf_in19.inv0.O buf_in19.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4234 VSS word2.buf_sel0.O word2.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4235 a_164100_3442# word3.byte1.tinv6.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4236 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4237 VDD word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4238 VDD a_108840_10088# a_108800_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4239 a_48180_2356# a_47970_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4240 VSS buf_sel7.inv0.O buf_sel7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4241 VDD a_105240_8628# word6.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4242 a_125910_9048# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4243 VDD word5.byte1.cgate0.nand0.B word5.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4244 VSS word5.byte1.tinv6.I a_164100_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4245 VDD buf_sel2.inv0.O buf_sel2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4246 a_101640_11764# a_101430_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4247 a_166050_11114# word8.byte1.dff_7.CLK a_165940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4248 a_141060_10088# a_140850_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4249 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4250 a_131700_7976# word6.byte1.cgate0.latch0.I0.ENB word6.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4251 VDD word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4252 VDD word3.byte1.cgate0.nand0.B word3.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4253 VSS word3.byte4.buf_RE0.O word3.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4254 a_116000_9598# a_115210_9548# a_115830_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4255 VSS a_65020_6412# a_64020_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4256 VDD word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4257 word8.byte3.dff_6.O word8.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4258 word8.gt_re3.I word8.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4259 word6.byte2.cgate0.nand0.A word6.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4260 VDD a_24420_6578# a_25980_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4261 a_112120_1090# a_110280_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4262 a_21820_7928# a_22150_8768# a_22050_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4263 VSS word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4264 buf_in28.inv1.O buf_in28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4265 VSS a_60420_4840# a_61980_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4266 a_124680_7976# word6.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4267 a_54220_6412# a_54550_6412# a_54450_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4268 VSS a_65020_3276# a_64020_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4269 VDD a_24420_3442# a_25980_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4270 Do22_buf buf_out23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4271 a_165100_6412# word5.byte1.dff_7.CLK a_165330_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4272 VSS word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4273 word6.byte3.cgate0.nand0.A word6.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4274 a_3820_140# word1.byte4.cgate0.inv1.O a_4050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4275 a_151260_190# word1.byte1.dff_7.CLK a_150700_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4276 word1.byte4.dff_6.O word1.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4277 VSS buf_in22.inv0.O buf_in22.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4278 a_42420_9714# word7.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4279 a_54220_3276# a_54550_3276# a_54450_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4280 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4281 VDD a_15780_680# word1.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4282 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4283 VSS CLK word2.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4284 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4285 VSS a_58980_680# a_58940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4286 a_165100_3276# word3.byte1.dff_7.CLK a_165330_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4287 a_147660_5912# word4.byte1.dff_7.CLK a_147100_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4288 a_128280_5796# word4.byte2.tinv7.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4289 VSS a_160500_9714# a_162060_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4290 a_47970_4842# word4.byte3.cgate0.inv1.O a_47860_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4291 a_140130_5912# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4292 a_50950_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4293 word4.byte3.dff_5.O word4.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4294 VDD word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4295 a_104080_4792# word4.byte2.dff_7.CLK a_104310_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4296 a_75360_10500# word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4297 a_161830_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4298 VSS a_126840_8628# word6.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4299 VDD a_62580_11764# word8.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4300 a_550_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4301 VDD word4.byte1.tinv3.I a_153300_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4302 VDD a_116040_10088# word7.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4303 a_50950_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4304 VDD buf_sel8.inv0.O buf_sel8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4305 a_158130_9048# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4306 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4307 a_104080_1656# word2.byte2.dff_7.CLK a_104310_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4308 a_19060_12184# a_17220_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4309 a_161830_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4310 a_48140_5912# a_47350_5632# a_47970_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4311 word6.byte4.dff_4.O word6.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4312 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4313 a_110280_4840# buf_out14.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4314 a_47250_4842# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4315 VDD a_142500_306# a_144060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4316 a_22150_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4317 a_53220_11112# buf_out21.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4318 VSS a_166260_680# word1.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4319 VDD word2.byte1.tinv3.I a_153300_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4320 VSS word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4321 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4322 a_112440_680# a_112230_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4323 VDD a_155460_5492# a_155420_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4324 a_100810_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4325 a_110280_1704# buf_out14.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4326 a_47250_1706# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4327 buf_out16.inv1.O buf_out16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4328 VSS word6.byte4.dff_0.O_bar a_2820_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4329 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4330 VDD word6.byte3.dff_0.O_bar a_42420_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4331 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4332 a_148220_9598# a_147430_9548# a_148050_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4333 VSS buf_out11.inv0.O buf_out11.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4334 a_28020_10500# buf_out25.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4335 VDD a_155460_2356# a_155420_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4336 a_100810_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4337 Do6_buf buf_out7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4338 Do27_buf buf_out28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4339 a_144340_7978# a_142500_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4340 word4.byte4.dff_1.O word4.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4341 a_55340_10498# word7.byte3.cgate0.inv1.O a_55170_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4342 VDD a_44580_8628# a_44540_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4343 a_118480_140# word1.byte2.dff_7.CLK a_118710_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4344 VSS word4.byte1.inv_and.O a_131700_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4345 VSS Di30 buf_in31.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4346 buf_in17.inv0.O Di16 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4347 a_15460_2776# a_13620_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4348 a_144060_7362# a_143830_6412# a_143500_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4349 word6.byte1.nand.B word6.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4350 a_44370_6462# a_43750_6412# a_44260_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4351 VDD a_111280_140# a_110280_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4352 a_147660_12184# word8.byte1.dff_7.CLK a_147100_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4353 VSS a_39720_7978# a_40380_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4354 VDD buf_out22.inv0.O Do21_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4355 a_107910_11114# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4356 a_151820_11114# word8.byte1.dff_7.CLK a_151650_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4357 VDD word5.byte1.cgate0.nand0.B word5.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4358 word2.byte4.dff_1.O word2.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4359 VSS a_1380_11764# word8.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4360 word5.byte3.dff_4.O word5.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4361 word4.byte1.dff_5.O word4.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4362 word6.byte3.tinv7.O word6.byte3.tinv1.EN a_46020_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4363 a_144060_4226# a_143830_3276# a_143500_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4364 word4.byte2.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B a_93540_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4365 a_154860_2776# word2.byte1.dff_7.CLK a_154300_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4366 a_44370_3326# a_43750_3276# a_44260_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4367 word5.byte1.tinv7.O buf_out7.inv0.I a_146100_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4368 VSS buf_sel2.inv0.O buf_sel2.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4369 word8.byte1.cgate0.inv1.I word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4370 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4371 a_2820_6578# word5.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4372 a_108240_190# word1.byte2.dff_7.CLK a_107680_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4373 a_17220_306# word1.byte4.tinv4.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4374 a_15780_2356# a_15570_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4375 word2.byte1.dff_5.O word2.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4376 VDD word3.byte1.cgate0.nand0.B word3.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4377 word3.byte3.dff_4.O word3.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4378 a_39180_5796# buf_we1.inv1.O word4.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4379 VDD word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4380 word6.byte2.dff_1.O word6.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4381 word3.byte1.tinv7.O buf_out7.inv0.I a_146100_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4382 a_119040_7978# a_118810_8768# a_118480_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4383 a_103080_3442# word3.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4384 a_95160_3442# word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4385 a_140130_12184# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4386 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4387 VSS word7.byte4.buf_RE0.O word7.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4388 a_150930_6462# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4389 VDD word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4390 a_19380_6952# a_19170_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4391 VSS word5.byte3.inv_and.O a_75720_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4392 a_55340_2776# a_54550_2496# a_55170_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4393 buf_in12.inv1.O buf_in12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4394 a_106680_11112# word8.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4395 a_159060_11764# a_158850_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4396 VDD word4.byte3.cgate0.nand0.A a_75360_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4397 a_17220_306# word1.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4398 a_139900_11064# word8.byte1.dff_7.CLK a_140130_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4399 a_26540_9048# a_25750_8768# a_26370_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4400 a_150930_3326# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4401 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4402 a_19380_3816# a_19170_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4403 a_166260_5492# a_166050_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4404 buf_in3.inv1.O buf_in3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4405 VDD a_21820_7928# a_20820_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4406 a_65350_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4407 VDD a_124680_11112# a_126240_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4408 VSS a_159060_11764# a_159020_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4409 a_58940_6462# a_58150_6412# a_58770_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4410 a_108010_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4411 VDD word2.byte3.cgate0.nand0.A a_75360_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4412 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.latch0.I0.O a_131700_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4413 a_10020_4840# word4.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4414 buf_in6.inv1.O buf_in6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4415 a_165940_9048# a_164100_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4416 a_8540_1090# word1.byte4.cgate0.inv1.O a_8370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4417 word2.byte1.tinv7.O word2.byte1.tinv6.EN a_164100_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4418 VDD word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4419 VSS word2.byte2.tinv2.I a_110280_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4420 a_58940_3326# a_58150_3276# a_58770_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4421 a_22150_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4422 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4423 VSS a_139800_11114# a_140460_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4424 a_165430_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4425 VDD buf_in18.inv0.O buf_in18.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4426 a_164100_4840# word4.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4427 buf_in30.inv1.O buf_in30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4428 a_126630_11114# word8.byte2.dff_7.CLK a_126520_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4429 VSS word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4430 a_101640_10088# a_101430_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4431 VSS word7.byte1.tinv0.I a_142500_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4432 VSS word1.byte4.buf_RE0.O word1.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4433 a_108800_4842# word4.byte2.dff_7.CLK a_108630_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4434 word8.byte1.tinv7.O buf_out7.inv0.I a_146100_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4435 VDD word7.byte2.buf_RE1.I word7.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4436 a_162620_7978# word6.byte1.dff_7.CLK a_162450_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4437 a_22050_1090# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4438 VSS a_111280_1656# a_110280_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4439 VDD a_26580_5492# word4.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4440 a_51460_6462# a_49620_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4441 VSS a_161500_140# a_160500_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4442 word4.byte3.tinv7.O word4.byte3.tinv3.EN a_53220_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4443 VSS word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4444 VSS word7.byte2.inv_and.O a_92280_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4445 VDD buf_sel3.inv0.O buf_sel3.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4446 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4447 a_108800_1706# word2.byte2.dff_7.CLK a_108630_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4448 a_1060_1090# a_120_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4449 VDD a_26580_2356# word2.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4450 a_156900_7976# buf_out4.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4451 a_56820_6578# word5.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4452 a_147430_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4453 a_51460_3326# a_49620_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4454 VSS a_151860_6952# word5.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4455 a_13620_6578# buf_out29.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4456 a_51780_6952# a_51570_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4457 VSS a_58980_10088# word7.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4458 a_36120_6578# word5.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4459 a_56820_3442# word3.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4460 a_162660_6952# a_162450_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4461 VSS a_151860_3816# word3.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4462 a_47020_7928# a_47350_8768# a_47250_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4463 word3.byte4.tinv7.O word3.byte4.tinv6.EN a_24420_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4464 a_13620_3442# buf_out29.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4465 a_51780_3816# a_51570_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4466 word6.byte3.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4467 a_1380_8628# a_1170_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4468 VSS word6.byte1.tinv2.I a_149700_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4469 a_162660_3816# a_162450_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4470 VSS a_141060_11764# word8.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4471 VSS word8.byte2.tinv2.I a_110280_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4472 VSS a_166260_11764# word8.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4473 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4474 a_106680_7976# word6.byte2.tinv1.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4475 a_18450_6462# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4476 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4477 a_164100_9714# word7.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4478 a_101640_5492# a_101430_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4479 VSS buf_in2.inv0.O buf_in2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4480 VDD a_42420_7976# a_43980_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4481 a_43750_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4482 VDD buf_out3.inv0.I buf_out3.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X4483 VDD a_62580_10088# word7.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4484 a_18450_3326# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4485 a_165330_5912# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4486 VSS word6.byte3.buf_RE0.O word6.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4487 a_101640_2356# a_101430_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4488 a_61980_1090# a_61750_140# a_61420_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4489 VSS dec8.and4_6.nand0.OUT buf_sel7.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4490 VDD word8.byte2.tinv6.I a_124680_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4491 a_22150_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4492 VSS a_113880_6578# a_115440_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4493 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4494 VDD buf_we3.inv0.O buf_we3.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4495 a_131700_1092# word1.byte1.cgate0.latch0.I0.ENB word1.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4496 VSS a_15780_10088# a_15740_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4497 a_149700_6578# word5.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4498 VSS a_113880_3442# a_115440_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4499 VDD word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4500 a_54780_11114# a_54550_11904# a_54220_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4501 a_149700_11112# buf_out6.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4502 a_124680_306# word1.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4503 word7.byte3.tinv7.O word7.byte3.tinv6.EN a_64020_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4504 VSS word5.byte2.buf_RE1.I word5.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4505 word5.byte2.tinv7.O word5.byte2.tinv1.EN a_106680_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4506 VSS a_108840_5492# a_108800_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4507 word1.byte2.cgate0.nand0.A word1.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4508 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4509 buf_sel5.inv1.O buf_sel5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4510 VSS a_118480_140# a_117480_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4511 VDD word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4512 VSS a_50620_6412# a_49620_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4513 VSS a_1380_2356# a_1340_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4514 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4515 VDD word6.byte3.tinv7.I a_67620_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4516 VDD a_10020_6578# a_11580_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4517 VDD word8.buf_sel0.O word8.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4518 VDD a_161500_6412# a_160500_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4519 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4520 a_116040_680# a_115830_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4521 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4522 VSS a_8580_680# a_8540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4523 a_7650_7362# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4524 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4525 VSS a_50620_3276# a_49620_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4526 word1.byte2.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4527 buf_re.inv1.O buf_re.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4528 word8.byte4.tinv7.O word8.byte4.tinv7.EN a_28020_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4529 VSS a_4980_6952# a_4940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4530 VDD a_10020_3442# a_11580_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4531 a_112400_11114# word8.byte2.dff_7.CLK a_112230_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4532 a_107910_10498# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4533 a_151820_10498# word7.byte1.dff_7.CLK a_151650_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4534 a_58380_6462# word5.byte3.cgate0.inv1.O a_57820_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4535 VDD a_161500_3276# a_160500_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4536 VSS buf_out27.inv0.O Do26_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4537 word7.byte4.dff_5.O word7.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4538 VSS buf_in8.inv0.O buf_in8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4539 a_7650_4226# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4540 VSS buf_out21.inv0.O Do20_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4541 VSS a_64020_7976# a_65580_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4542 VSS a_4980_3816# a_4940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4543 a_58380_3326# word3.byte3.cgate0.inv1.O a_57820_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4544 a_113880_4840# word4.byte2.tinv3.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4545 word4.byte2.dff_3.O word4.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4546 VDD buf_out2.inv0.O Do1_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4547 a_7980_7978# a_7750_8768# a_7420_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4548 VSS a_166260_5492# word4.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4549 VDD a_40980_11764# a_40940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4550 VDD a_66180_11764# a_66140_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4551 VDD word5.byte2.tinv4.I a_117480_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4552 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4553 VSS word2.byte4.cgate0.latch0.I0.O word2.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4554 a_111610_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4555 a_75720_5796# word4.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4556 word5.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4557 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4558 a_162060_7978# a_161830_8768# a_161500_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4559 a_62370_7978# a_61750_8768# a_62260_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4560 a_143730_9048# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4561 word7.byte1.cgate0.inv1.I word7.byte1.cgate0.nand0.A a_134580_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4562 a_128280_3442# word3.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4563 VDD word3.byte2.tinv4.I a_117480_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4564 VDD a_157900_4792# a_156900_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4565 VDD word4.byte1.buf_RE1.I word4.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4566 a_159060_10088# a_158850_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4567 VSS word4.byte1.cgate0.nand0.B a_33420_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4568 a_139900_9548# word7.byte1.dff_7.CLK a_140130_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4569 word5.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4570 VDD word5.byte1.cgate0.nand0.B word5.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4571 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4572 VSS word1.byte1.tinv2.I a_149700_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4573 VDD a_105240_6952# a_105200_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4574 a_101430_7978# word6.byte2.dff_7.CLK a_101320_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4575 word3.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4576 word3.byte2.nand.OUT buf_we3.inv1.O a_90120_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4577 word3.byte3.inv_and.O word3.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4578 VSS a_11020_4792# a_10020_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4579 VDD a_124680_9714# a_126240_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4580 VDD word5.byte4.inv_and.O a_36120_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4581 VDD word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4582 word6.byte1.tinv7.O buf_out6.inv0.I a_149700_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4583 VDD a_157900_1656# a_156900_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4584 VDD word1.byte3.dff_0.O_bar a_42420_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4585 VDD word2.byte1.buf_RE1.I word2.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4586 VDD word3.byte1.cgate0.nand0.B word3.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4587 word3.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4588 VDD a_220_4792# a_120_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4589 VSS word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4590 VDD a_105240_3816# a_105200_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4591 a_158230_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4592 a_60420_11112# word8.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4593 VDD word3.byte4.inv_and.O a_36120_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4594 VSS buf_in9.inv0.O buf_in9.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4595 a_28020_7976# word6.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4596 VSS word5.byte4.tinv4.I a_17220_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4597 VDD a_220_1656# a_120_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4598 a_158230_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4599 buf_in28.inv1.O buf_in28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4600 a_4980_11764# a_4770_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4601 a_122640_9598# word7.byte2.dff_7.CLK a_122080_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4602 VSS a_161500_7928# a_160500_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4603 a_142500_7976# word6.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4604 a_148260_8628# a_148050_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4605 buf_in5.inv0.O Di4 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4606 VSS buf_in17.inv0.O buf_in17.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4607 word8.byte2.tinv7.O buf_out15.inv0.I a_106680_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4608 a_47350_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4609 a_155250_190# word1.byte1.dff_7.CLK a_155140_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4610 VSS word6.byte2.buf_RE1.I word6.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4611 a_92280_8932# word6.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4612 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4613 VSS word8.byte1.tinv7.I a_167700_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4614 VSS a_14620_140# a_13620_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4615 VDD buf_in20.inv0.O buf_in20.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4616 word5.byte3.dff_0.O word5.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4617 a_115110_1090# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4618 VSS word7.byte1.tinv7.I a_167700_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4619 a_44260_9048# a_42420_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4620 VSS word3.byte4.tinv1.I a_6420_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4621 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.latch0.I0.O a_132960_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4622 word2.byte2.dff_5.O word2.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4623 a_124680_9714# word7.byte2.tinv6.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4624 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4625 a_18220_6412# word5.byte4.cgate0.inv1.O a_18450_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4626 a_104640_1090# a_104410_140# a_104080_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4627 word3.byte3.dff_0.O word3.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4628 VSS a_39820_1656# a_39720_1706# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4629 a_74100_13636# dec8.and4_5.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4630 a_132960_306# word1.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4631 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4632 VSS a_144660_8628# word6.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4633 word8.byte2.dff_5.O word8.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4634 a_75360_9714# word7.byte1.cgate0.nand0.B word7.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4635 VSS word3.buf_ck1.I word3.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4636 a_54220_4792# a_54550_5632# a_54450_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4637 buf_sel5.inv1.O buf_sel5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4638 a_14950_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4639 a_46020_11112# buf_out23.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4640 a_44580_8628# a_44370_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4641 word1.byte1.tinv7.O word1.byte1.tinv1.EN a_146100_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4642 word5.byte1.inv_and.O word5.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4643 a_18220_3276# word3.byte4.cgate0.inv1.O a_18450_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4644 VSS a_13620_9714# a_15180_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4645 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4646 VSS word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4647 VSS a_165100_9548# a_164100_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4648 a_40940_2776# a_40150_2496# a_40770_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4649 VSS a_101640_11764# word8.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4650 a_49620_3442# word3.byte3.tinv2.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4651 a_14950_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4652 a_11020_7928# word6.byte4.cgate0.inv1.O a_11250_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4653 a_154300_9548# a_154630_9548# a_154530_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4654 a_112400_6462# a_111610_6412# a_112230_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4655 a_50950_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4656 a_22660_11114# a_20820_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4657 a_60420_7976# word6.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4658 VSS a_148260_2356# a_148220_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4659 a_132960_8932# word6.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4660 a_14950_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4661 VDD buf_out11.inv0.I buf_out11.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X4662 VSS word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4663 a_112400_3326# a_111610_3276# a_112230_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4664 VDD a_147100_140# a_146100_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4665 a_126840_5492# a_126630_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4666 VSS buf_out2.inv0.I buf_out2.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X4667 VSS a_2820_6578# a_4380_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4668 word7.byte4.inv_and.O word7.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4669 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4670 VSS word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4671 VSS word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4672 VSS a_39820_140# a_39720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4673 Do30_buf buf_out31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4674 VDD buf_in4.inv0.O buf_in4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4675 a_126840_2356# a_126630_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4676 VSS a_106680_7976# a_108240_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4677 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4678 VSS a_2820_3442# a_4380_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4679 a_148050_4842# a_147430_5632# a_147940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4680 a_110280_11112# buf_out14.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4681 VDD word7.byte3.tinv6.I a_64020_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4682 a_17220_11112# word8.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4683 a_54780_10498# a_54550_9548# a_54220_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4684 VDD a_116040_8628# word6.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4685 a_56820_1704# word2.byte3.tinv4.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4686 VSS word6.byte4.tinv2.I a_10020_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4687 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4688 a_780_9598# word7.byte4.cgate0.inv1.O a_220_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4689 a_156900_306# buf_out4.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4690 a_147330_7978# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4691 a_110280_6578# word5.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4692 a_148050_1706# a_147430_2496# a_147940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4693 a_158130_12184# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4694 word4.byte4.tinv7.O buf_out31.inv0.I a_6420_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4695 buf_sel7.inv1.O buf_sel7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4696 VSS a_56820_306# a_58380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4697 a_110280_3442# word3.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4698 a_61420_1656# a_61750_2496# a_61650_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4699 word8.byte4.dff_6.O word8.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4700 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4701 word4.byte4.dff_3.O word4.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4702 word8.byte3.dff_2.O word8.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4703 word5.byte1.dff_4.O word5.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4704 a_65250_190# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4705 word2.byte4.tinv7.O buf_out31.inv0.I a_6420_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4706 VSS word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4707 word1.byte3.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4708 a_122920_1090# a_121080_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4709 VDD word4.byte3.buf_RE0.O word4.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4710 a_157900_11064# word8.byte1.dff_7.CLK a_158130_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4711 a_112400_10498# word7.byte2.dff_7.CLK a_112230_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4712 VDD a_139800_4842# a_140460_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4713 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4714 a_22980_11764# a_22770_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4715 a_158230_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4716 word3.byte4.tinv7.O word3.byte4.tinv2.EN a_10020_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4717 word2.byte4.dff_3.O word2.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4718 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4719 word3.byte1.dff_4.O word3.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4720 VDD word2.byte3.buf_RE0.O word2.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4721 VDD a_139800_1706# a_140460_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4722 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4723 VDD a_40980_10088# a_40940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4724 a_117480_306# word1.byte2.tinv4.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4725 word7.byte3.dff_1.O word7.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4726 VDD a_66180_10088# a_66140_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4727 VSS buf_out8.inv0.O Do7_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4728 VSS buf_in20.inv0.O buf_in20.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4729 a_56820_306# word1.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4730 a_10020_11112# word8.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4731 VSS a_156900_11112# a_158460_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4732 VDD buf_we2.inv0.O buf_we2.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4733 buf_in1.inv0.O Di0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4734 a_150930_5912# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4735 VDD a_162660_11764# a_162620_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4736 VSS a_147100_1656# a_146100_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4737 a_19380_5492# a_19170_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4738 buf_in22.inv1.O buf_in22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4739 a_15570_190# a_14950_140# a_15460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4740 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4741 a_90120_2660# word2.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4742 a_160500_9714# word7.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4743 word6.byte4.dff_0.O word6.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4744 VSS a_40980_680# a_40940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4745 a_119320_6462# a_117480_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4746 word1.byte4.dff_7.O word1.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4747 VDD a_148260_8628# word6.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4748 word2.byte4.tinv7.O word2.byte4.tinv4.EN a_17220_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4749 a_58940_5912# a_58150_5632# a_58770_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4750 a_58050_4842# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4751 VDD a_153300_306# a_154860_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4752 a_121080_4840# buf_out11.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4753 a_126630_7978# word6.byte2.dff_7.CLK a_126520_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4754 a_18550_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4755 a_119320_3326# a_117480_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4756 VDD word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4757 a_115440_4842# a_115210_5632# a_114880_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4758 a_17220_4840# word4.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4759 a_4050_190# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4760 VDD word1.byte3.tinv7.I a_67620_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4761 VDD word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4762 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4763 VSS word8.buf_ck1.I word8.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4764 VDD word6.byte2.tinv5.I a_121080_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4765 a_58050_1706# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4766 a_121080_1704# buf_out11.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4767 a_4980_10088# a_4770_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4768 word3.byte3.cgate0.inv1.I word3.byte3.cgate0.nand0.A a_73020_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4769 word4.gt_re3.I word4.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4770 a_15740_7978# word6.byte4.cgate0.inv1.O a_15570_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4771 VDD word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4772 a_40380_2776# word2.byte3.cgate0.inv1.O a_39820_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4773 VDD word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4774 a_115440_1706# a_115210_2496# a_114880_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4775 a_159020_9598# a_158230_9548# a_158850_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4776 a_4150_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4777 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4778 VDD word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4779 a_15460_7362# a_13620_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4780 a_155140_1090# a_153300_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4781 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4782 VDD a_55380_680# a_55340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4783 a_11580_9048# word6.byte4.cgate0.inv1.O a_11020_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4784 VDD a_123240_8628# a_123200_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4785 word2.gt_re3.I word2.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4786 VDD buf_in13.inv0.O buf_in13.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4787 VDD word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4788 VSS a_159060_11764# word8.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4789 VDD a_122080_7928# a_121080_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4790 a_51460_5912# a_49620_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4791 VSS word8.byte2.tinv7.I a_128280_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4792 a_43980_6462# word5.byte3.cgate0.inv1.O a_43420_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4793 VDD word8.byte2.cgate0.nand0.A word8.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4794 a_167700_8932# word6.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4795 a_156900_9714# word7.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4796 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4797 a_15460_4226# a_13620_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4798 VSS buf_in4.inv0.O buf_in4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4799 word7.byte4.tinv7.O buf_out27.inv0.I a_20820_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4800 a_7750_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4801 a_6420_1704# word2.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4802 a_154860_7362# a_154630_6412# a_154300_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4803 VSS buf_in25.inv0.O buf_in25.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4804 word6.byte2.tinv7.O word6.byte2.tinv6.EN a_124680_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4805 a_15780_6952# a_15570_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4806 a_43980_3326# word3.byte3.cgate0.inv1.O a_43420_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4807 VSS word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4808 VSS a_151860_5492# word4.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4809 a_153300_11112# word8.byte1.tinv3.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4810 a_4940_4842# word4.byte4.cgate0.inv1.O a_4770_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4811 a_154860_4226# a_154630_3276# a_154300_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4812 a_7750_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4813 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4814 a_51780_5492# a_51570_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4815 a_14950_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4816 a_15780_3816# a_15570_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4817 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4818 word1.gt_re0.OUT buf_sel1.inv1.O a_82020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4819 a_48140_190# a_47350_140# a_47970_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4820 a_4940_1706# word2.byte4.cgate0.inv1.O a_4770_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4821 a_147100_4792# word4.byte1.dff_7.CLK a_147330_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4822 a_55340_7362# word5.byte3.cgate0.inv1.O a_55170_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4823 VDD EN dec8.and4_7.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4824 word2.byte3.tinv7.O word2.byte3.tinv2.EN a_49620_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4825 a_113880_3442# word3.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4826 a_167700_11112# buf_out1.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4827 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4828 word1.byte1.tinv7.O buf_out6.inv0.I a_149700_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4829 VDD word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4830 a_151860_10088# a_151650_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4831 a_147100_1656# word2.byte1.dff_7.CLK a_147330_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4832 VSS word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4833 a_55340_4226# word3.byte3.cgate0.inv1.O a_55170_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4834 a_18450_5912# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4835 a_153300_4840# buf_out5.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4836 word8.byte2.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B a_93540_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4837 a_22660_10498# a_20820_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4838 a_108010_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4839 a_105200_9048# a_104410_8768# a_105030_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4840 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4841 a_28020_1092# word1.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4842 a_143830_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4843 VSS a_118480_6412# a_117480_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4844 a_143500_140# a_143830_140# a_143730_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4845 VSS a_55380_6952# word5.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4846 a_153300_1704# buf_out5.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4847 VSS buf_out10.inv0.I buf_out10.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X4848 a_108010_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4849 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4850 a_118810_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4851 VDD word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4852 a_65250_11114# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4853 a_143830_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4854 a_2820_7976# word6.byte4.tinv0.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4855 VSS a_113880_4840# a_115440_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4856 Do5_buf buf_out6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4857 VSS a_118480_3276# a_117480_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4858 a_42420_7976# buf_out24.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4859 VSS a_55380_3816# word3.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4860 VDD a_4980_8628# word6.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4861 VSS buf_out23.inv0.O Do22_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4862 VSS buf_in3.inv0.O buf_in3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4863 VDD a_14620_6412# a_13620_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4864 a_100710_1090# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4865 VDD a_58980_11764# a_58940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4866 VDD word7.byte1.tinv5.I a_160500_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4867 a_131700_5796# word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4868 dec8.and4_0.nand1.OUT dec8.and4_3.nand1.A a_64560_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4869 VDD a_14620_3276# a_13620_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4870 buf_in18.inv1.O buf_in18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4871 word7.byte4.dff_6.O word7.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4872 word7.byte3.dff_2.O word7.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4873 word4.byte2.cgate0.nand0.A word4.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4874 buf_sel8.inv1.O buf_sel8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4875 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4876 a_157900_9548# word7.byte1.dff_7.CLK a_158130_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4877 word5.byte4.tinv7.O word5.byte4.tinv0.EN a_2820_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4878 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4879 a_115440_190# word1.byte2.dff_7.CLK a_114880_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4880 a_26370_4842# a_25750_5632# a_26260_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4881 VSS a_4980_5492# a_4940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4882 VDD a_64020_11112# a_65580_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4883 word6.byte1.dff_2.O word6.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4884 VSS a_12180_6952# a_12140_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4885 a_24420_306# word1.byte4.tinv6.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4886 a_146100_3442# word3.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4887 a_58380_5912# word4.byte3.cgate0.inv1.O a_57820_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4888 VSS a_150700_9548# a_149700_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4889 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4890 word8.byte1.dff_1.O word8.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X4891 VDD word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4892 CLK buf_ck.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4893 a_125680_7928# a_126010_8768# a_125910_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X4894 a_19060_9598# a_17220_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4895 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4896 a_26370_1706# a_25750_2496# a_26260_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4897 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4898 a_25650_2776# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4899 VDD a_164100_4840# a_165660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4900 a_60420_306# word1.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4901 VSS a_12180_3816# a_12140_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4902 a_144660_11764# a_144450_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4903 VSS word3.byte4.cgate0.nand0.A a_35760_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4904 a_151650_6462# word5.byte1.dff_7.CLK a_151540_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4905 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4906 VSS word5.byte1.cgate0.nand0.B word5.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4907 a_450_1090# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X4908 VDD word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4909 VSS buf_out16.inv0.O buf_out16.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4910 VSS a_119640_10088# word7.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4911 a_15180_7978# a_14950_8768# a_14620_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4912 VDD word4.byte3.tinv6.I a_64020_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4913 VDD word6.byte4.cgate0.nand0.A word6.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4914 a_158460_9598# word7.byte1.dff_7.CLK a_157900_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4915 a_58770_9598# word7.byte3.cgate0.inv1.O a_58660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4916 VDD a_164100_1704# a_165660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4917 buf_in9.inv0.O buf_in9.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4918 a_65970_11114# word8.byte3.cgate0.inv1.O a_65860_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4919 a_151650_3326# word3.byte1.dff_7.CLK a_151540_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4920 a_3820_11064# word8.byte4.cgate0.inv1.O a_4050_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X4921 VDD a_123240_11764# a_123200_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4922 VDD a_162660_10088# a_162620_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4923 a_122410_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X4924 VDD word2.byte3.tinv6.I a_64020_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4925 a_112440_5492# a_112230_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4926 VSS a_121080_1704# a_122640_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4927 VDD a_53220_7976# a_54780_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4928 VDD a_66180_5492# a_66140_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4929 VSS word2.byte1.tinv3.I a_153300_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4930 a_8260_6462# a_6420_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4931 VDD buf_out5.inv0.O Do4_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4932 a_112440_2356# a_112230_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4933 VDD a_101640_680# word1.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X4934 a_110280_1704# word2.byte2.tinv2.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4935 VSS a_6420_306# a_7980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4936 VDD a_66180_2356# a_66140_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4937 Do21_buf buf_out22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4938 a_4380_4842# a_4150_5632# a_3820_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4939 VSS word6.byte1.cgate0.nand0.B word6.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4940 a_8260_3326# a_6420_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4941 VSS a_2820_11112# a_4380_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X4942 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4943 a_66900_13636# dec8.and4_1.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4944 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4945 VSS a_14620_7928# a_13620_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4946 a_8580_6952# a_8370_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4947 a_142500_9714# word7.byte1.tinv0.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X4948 VDD a_1380_6952# a_1340_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4949 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4950 VDD word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4951 a_4380_1706# a_4150_2496# a_3820_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X4952 VSS word4.byte3.dff_0.O_bar a_42420_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4953 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4954 VSS a_15780_680# word1.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4955 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4956 a_92280_9714# word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4957 VDD word5.byte2.buf_RE1.I word5.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4958 a_8580_3816# a_8370_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X4959 VDD word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4960 VSS word8.gt_re1.O word8.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4961 VDD buf_sel6.inv0.I buf_sel6.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4962 VDD a_1380_3816# a_1340_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X4963 VSS word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4964 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4965 word5.byte3.tinv7.O buf_out20.inv0.I a_56820_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4966 a_65580_2776# word2.byte3.cgate0.inv1.O a_65020_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4967 VDD word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4968 VDD word3.byte2.buf_RE1.I word3.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4969 a_117480_9714# word7.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4970 a_6420_306# word1.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4971 VSS buf_in12.inv0.O buf_in12.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4972 word3.byte3.tinv7.O buf_out20.inv0.I a_56820_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4973 word5.byte4.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4974 VSS a_100480_140# a_100380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X4975 VDD a_43420_4792# a_42420_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4976 a_24420_4840# word4.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4977 word8.gt_re0.OUT buf_sel8.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4978 a_61650_6462# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4979 word7.byte1.tinv7.O buf_out8.inv0.I a_142500_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4980 a_11580_190# word1.byte4.cgate0.inv1.O a_11020_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4981 VSS buf_in8.inv0.O buf_in8.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X4982 VSS a_18220_9548# a_17220_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X4983 VDD a_43420_1656# a_42420_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X4984 a_24420_1704# word2.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4985 a_144660_5492# a_144450_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4986 VDD buf_in29.inv0.O buf_in29.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4987 a_101320_2776# a_100380_1706# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4988 a_61650_3326# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X4989 VDD buf_in23.inv0.O buf_in23.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X4990 a_2820_9714# word7.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X4991 VDD word7.byte3.tinv4.I a_56820_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4992 buf_in18.inv1.O buf_in18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X4993 a_103080_11112# buf_out16.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X4994 a_128280_11112# buf_out9.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4995 a_144660_2356# a_144450_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X4996 word7.byte1.cgate0.nand0.A word7.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4997 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X4998 a_112400_5912# a_111610_5632# a_112230_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X4999 a_104920_6462# a_103080_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5000 a_111510_4842# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5001 VSS word2.byte3.cgate0.nand0.A a_75360_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5002 word1.byte4.cgate0.inv1.I word1.byte4.cgate0.nand0.A a_33420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5003 VSS a_120_1706# a_780_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5004 word7.gt_re1.O word7.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5005 VSS a_7420_6412# a_6420_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5006 a_158740_190# a_156900_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5007 VDD word1.byte2.tinv5.I a_121080_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5008 VSS a_21820_4792# a_20820_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5009 a_40380_12184# word8.byte3.cgate0.inv1.O a_39820_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5010 word7.byte2.cgate0.inv1.I word7.byte2.cgate0.nand0.A a_95160_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5011 a_111510_1706# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5012 a_104920_3326# a_103080_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5013 a_101040_4842# a_100810_5632# a_100480_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5014 a_149700_6578# word5.byte1.tinv2.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5015 buf_sel4.inv0.I dec8.and4_3.nand1.OUT a_70500_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5016 VSS a_2820_4840# a_4380_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5017 a_65250_10498# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5018 VSS a_48180_8628# word6.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5019 VSS a_7420_3276# a_6420_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5020 VSS word7.byte3.tinv3.I a_53220_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5021 VDD word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5022 a_106680_7976# word6.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5023 VSS word1.byte1.inv_and.O a_131700_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5024 a_101040_1706# a_100810_2496# a_100480_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5025 word7.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5026 a_21820_11064# a_22150_11904# a_22050_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5027 a_140740_1090# a_139800_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5028 a_161730_11114# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5029 VDD a_40980_680# a_40940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5030 VSS a_125680_140# a_124680_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5031 a_150700_6412# a_151030_6412# a_150930_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5032 a_159060_680# a_158850_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5033 VDD buf_out12.inv0.O buf_out12.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5034 a_67620_7976# buf_out17.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5035 a_58150_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5036 word8.byte2.cgate0.nand0.A word8.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5037 VDD a_58980_10088# a_58940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5038 a_126010_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5039 VDD word7.byte2.tinv5.I a_121080_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5040 word1.byte3.dff_7.O word1.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5041 a_150700_3276# a_151030_3276# a_150930_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5042 word5.byte2.dff_5.O word5.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5043 word6.byte2.tinv7.O word6.byte2.tinv2.EN a_110280_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5044 a_51780_11764# a_51570_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5045 VSS word8.byte1.cgate0.nand0.B a_134580_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5046 VDD a_39820_6412# a_39720_6462# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5047 a_125910_1090# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5048 a_39820_9548# a_40150_9548# a_40050_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5049 a_156900_4840# word4.byte1.tinv4.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5050 word3.byte2.dff_5.O word3.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5051 word4.byte1.dff_4.O word4.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5052 VSS buf_in31.inv0.O buf_in31.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5053 buf_in17.inv1.O buf_in17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5054 VDD a_64020_9714# a_65580_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5055 VDD a_39820_3276# a_39720_3326# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5056 VDD buf_out32.inv0.O Do31_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5057 a_160500_11112# word8.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5058 a_40940_7362# word5.byte3.cgate0.inv1.O a_40770_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5059 word8.byte2.dff_1.O word8.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5060 word7.byte1.dff_1.O word7.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5061 VDD a_112440_5492# word4.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5062 a_450_11114# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5063 a_55380_8628# a_55170_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5064 a_117480_6578# buf_out12.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5065 VDD word8.byte4.tinv3.I a_13620_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5066 VSS a_100480_1656# a_100380_1706# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5067 a_40940_4226# word3.byte3.cgate0.inv1.O a_40770_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5068 word4.byte3.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5069 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5070 VDD a_112440_2356# word2.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5071 buf_sel1.inv1.O buf_sel1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5072 a_21820_140# word1.byte4.cgate0.inv1.O a_22050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5073 VSS word8.byte2.buf_RE1.I word8.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5074 VDD word5.buf_ck1.I word5.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5075 VDD a_148260_6952# a_148220_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5076 a_144450_7978# word6.byte1.dff_7.CLK a_144340_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5077 a_117480_3442# buf_out12.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5078 VDD word4.byte1.buf_RE1.I word4.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5079 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5080 a_3820_9548# word7.byte4.cgate0.inv1.O a_4050_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5081 VDD a_123240_10088# a_123200_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5082 VDD word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5083 buf_in15.inv0.O buf_in15.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5084 a_13620_9714# word7.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5085 VSS a_40980_6952# word5.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5086 a_108240_2776# word2.byte2.dff_7.CLK a_107680_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5087 VDD a_148260_3816# a_148220_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5088 VDD word3.buf_ck1.I word3.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5089 word4.byte1.nand.B word4.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5090 VSS word5.byte3.tinv5.I a_60420_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5091 a_42420_306# buf_out24.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5092 VDD word2.byte1.buf_RE1.I word2.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5093 VDD buf_we4.inv0.O buf_we4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5094 word1.byte4.dff_1.O word1.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5095 VDD a_157900_140# a_156900_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5096 VSS a_40980_3816# word3.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5097 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5098 VDD a_141060_8628# a_141020_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5099 a_123200_190# a_122410_140# a_123030_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5100 word2.byte1.nand.B word2.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5101 a_119320_5912# a_117480_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5102 VSS buf_re.inv0.O buf_re.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5103 word6.byte4.tinv7.O buf_out25.inv0.I a_28020_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5104 a_17220_6578# word5.byte4.tinv4.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5105 VDD a_120_11114# a_780_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5106 VSS word6.byte1.cgate0.nand0.B word6.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5107 VDD buf_in4.inv0.O buf_in4.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5108 a_146100_11112# word8.byte1.tinv1.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5109 VDD a_126840_680# word1.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5110 word6.byte1.tinv7.O word6.byte1.tinv0.EN a_142500_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5111 VSS word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5112 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5113 a_158130_1090# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5114 VSS word6.byte4.tinv5.I a_20820_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5115 a_162450_190# word1.byte1.dff_7.CLK a_162340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5116 VSS a_119640_10088# a_119600_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5117 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5118 Do18_buf buf_out19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5119 VSS a_40980_11764# word8.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5120 a_61420_6412# word5.byte3.cgate0.inv1.O a_61650_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5121 VSS a_21820_140# a_20820_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5122 word2.byte1.dff_6.O word2.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5123 VSS a_66180_11764# word8.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5124 a_167700_9714# word7.byte1.tinv7.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5125 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5126 VSS word4.byte3.tinv7.I a_67620_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5127 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5128 a_6420_3442# word3.byte4.tinv1.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5129 a_11970_4842# a_11350_5632# a_11860_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5130 buf_sel7.inv1.O buf_sel7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5131 a_115830_7978# a_115210_8768# a_115720_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5132 VDD word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5133 a_108630_190# word1.byte2.dff_7.CLK a_108520_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5134 a_131700_3442# word3.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5135 a_61420_3276# word3.byte3.cgate0.inv1.O a_61650_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5136 a_43980_5912# word4.byte3.cgate0.inv1.O a_43420_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5137 word4.byte4.dff_6.O word4.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5138 VDD buf_out17.inv0.O Do16_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5139 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5140 VDD word5.gt_re0.OUT word5.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5141 a_7750_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5142 VDD buf_sel3.inv0.I buf_sel3.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5143 a_111280_7928# a_111610_8768# a_111510_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5144 word1.gt_re3.I word1.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5145 a_75720_9714# word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5146 a_11970_1706# a_11350_2496# a_11860_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5147 VSS word3.buf_ck1.I word3.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5148 VDD word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5149 VDD word1.byte4.cgate0.nand0.A word1.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5150 word1.byte1.tinv7.O word1.byte1.tinv3.EN a_153300_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5151 VSS buf_out12.inv0.I buf_out12.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X5152 word2.byte4.dff_6.O word2.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5153 a_93540_3442# word3.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5154 VDD word3.gt_re0.OUT word3.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5155 VSS a_39720_190# a_40380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5156 a_12140_4842# word4.byte4.cgate0.inv1.O a_11970_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5157 a_58050_11114# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5158 a_155140_11114# a_153300_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5159 a_54450_9048# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5160 a_155420_6462# a_154630_6412# a_155250_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5161 VDD buf_in16.inv0.O buf_in16.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5162 a_49620_4840# word4.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5163 word7.byte2.dff_6.O word7.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5164 a_20820_6578# word5.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5165 VDD a_39720_190# a_40380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5166 VSS a_162660_8628# a_162620_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5167 a_140230_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5168 a_12140_1706# word2.byte4.cgate0.inv1.O a_11970_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5169 a_151540_4842# a_149700_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5170 VSS buf_in28.inv0.O buf_in28.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5171 a_155420_3326# a_154630_3276# a_155250_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5172 word6.byte3.tinv7.O buf_out19.inv0.I a_60420_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5173 a_49620_1704# word2.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5174 VDD a_51780_5492# a_51740_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5175 VDD buf_out23.inv0.I buf_out23.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X5176 a_58660_7978# a_56820_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5177 a_126520_2776# a_124680_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5178 VSS a_157900_1656# a_156900_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5179 VSS word2.byte1.buf_RE1.I word2.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5180 a_151540_1706# a_149700_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5181 a_155420_12184# a_154630_11904# a_155250_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5182 a_44540_9598# a_43750_9548# a_44370_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5183 word6.gt_re3.I word6.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5184 a_122640_11114# a_122410_11904# a_122080_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5185 a_42420_9714# buf_out24.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5186 VDD a_51780_2356# a_51740_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5187 buf_in22.inv1.O buf_in22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5188 word1.byte2.dff_1.O word1.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5189 word4.byte1.tinv7.O word4.byte1.tinv2.EN a_149700_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5190 VSS word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5191 a_56820_11112# word8.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5192 buf_we2.inv1.O buf_we2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5193 VDD a_159060_8628# word6.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5194 VSS a_55380_5492# word4.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5195 a_53220_7976# word6.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5196 a_58980_8628# a_58770_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5197 a_40380_7362# a_40150_6412# a_39820_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5198 a_153300_6578# word5.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5199 buf_sel6.inv0.I dec8.and4_5.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5200 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5201 a_4150_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5202 a_28020_5796# word4.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5203 a_162060_12184# word8.byte1.dff_7.CLK a_161500_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5204 a_1340_9048# a_550_8768# a_1170_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5205 a_26540_1090# word1.byte4.cgate0.inv1.O a_26370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5206 buf_sel8.inv1.O buf_sel8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5207 a_122920_12184# a_121080_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5208 a_122310_11114# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5209 a_161730_10498# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5210 VSS word1.buf_ck1.I word1.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5211 VSS word3.gt_re1.O word3.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5212 word7.byte2.inv_and.O word7.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5213 VDD a_12180_8628# word6.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5214 a_153300_3442# word3.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5215 a_40380_4226# a_40150_3276# a_39820_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5216 a_19170_1706# word2.byte4.cgate0.inv1.O a_19060_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5217 a_4150_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5218 word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.latch0.I0.O a_36120_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5219 VSS a_64020_306# a_65580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5220 VSS word3.byte4.buf_RE0.O word3.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5221 a_165940_1090# a_164100_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5222 VSS a_103080_11112# a_104640_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5223 a_129540_12068# word8.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5224 VSS word5.byte1.cgate0.nand0.B a_95160_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5225 a_51780_10088# a_51570_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5226 word6.byte4.nand.OUT word6.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5227 VSS a_156900_1704# a_158460_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5228 a_165430_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5229 VDD word7.byte4.buf_RE0.O word7.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5230 VSS buf_out25.inv0.O Do24_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5231 a_140230_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5232 VDD buf_out7.inv0.O Do6_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5233 VDD a_17220_4840# a_18780_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5234 VDD a_1380_5492# word4.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5235 VDD buf_out28.inv0.I buf_out28.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X5236 a_121080_11112# word8.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5237 VSS a_12180_5492# a_12140_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5238 word7.byte2.dff_1.O word7.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5239 a_62580_680# a_62370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5240 a_124680_306# word1.byte2.tinv6.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5241 a_65020_9548# a_65350_9548# a_65250_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5242 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5243 a_105240_2356# a_105030_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5244 a_450_10498# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5245 VSS buf_out31.inv0.O Do30_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5246 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5247 VSS word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5248 a_64020_306# word1.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5249 VDD a_17220_1704# a_18780_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5250 VDD a_1380_2356# word2.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5251 a_151650_4842# word4.byte1.dff_7.CLK a_151540_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5252 word8.byte4.cgate0.nand0.A word8.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5253 word7.buf_sel0.O buf_sel7.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X5254 buf_sel3.inv1.O buf_sel3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5255 VSS a_62580_2356# word2.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5256 a_61750_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5257 word7.byte1.tinv7.O word7.byte1.tinv5.EN a_160500_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5258 VSS word1.byte2.inv_and.O a_92280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5259 a_164100_4840# buf_out2.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5260 a_118810_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5261 a_47020_140# word1.byte3.cgate0.inv1.O a_47250_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5262 VDD word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5263 a_106680_306# word1.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5264 a_60420_4840# word4.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5265 VSS word8.byte3.tinv5.I a_60420_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5266 a_116000_9048# a_115210_8768# a_115830_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5267 a_114880_7928# word6.byte2.dff_7.CLK a_115110_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5268 VSS a_100380_9598# a_101040_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5269 VSS word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5270 word8.byte1.tinv7.O buf_out3.inv0.I a_160500_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5271 a_8260_5912# a_6420_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5272 VDD word6.byte1.tinv6.I a_164100_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5273 a_164100_1704# buf_out2.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5274 VDD word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5275 a_118810_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5276 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5277 a_67620_1092# buf_out17.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5278 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5279 VDD a_120_9598# a_780_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5280 VDD buf_in12.inv0.O buf_in12.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5281 a_106680_11112# word8.byte2.tinv1.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5282 a_43750_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5283 VDD word4.byte4.buf_RE0.O word4.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5284 a_111610_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5285 VDD a_166260_8628# a_166220_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5286 VDD word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5287 a_55170_6462# word5.byte3.cgate0.inv1.O a_55060_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5288 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5289 a_8580_5492# a_8370_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5290 VSS buf_in3.inv0.O buf_in3.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5291 VSS a_160500_7976# a_162060_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5292 word5.byte3.dff_7.O word5.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5293 a_1380_680# a_1170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5294 VDD buf_in10.inv0.I buf_in10.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5295 VDD word2.byte4.buf_RE0.O word2.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5296 VDD buf_we1.inv0.O buf_we1.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5297 a_55170_3326# word3.byte3.cgate0.inv1.O a_55060_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5298 VDD a_49620_4840# a_51180_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5299 word6.byte1.tinv7.O word6.byte1.tinv7.EN a_167700_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5300 a_4770_7978# a_4150_8768# a_4660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5301 VSS word6.byte2.tinv3.I a_113880_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5302 VSS a_101640_680# word1.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5303 VSS Di0 buf_in1.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5304 word7.byte4.cgate0.inv1.I word7.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5305 word2.byte4.tinv7.O word2.byte4.tinv1.EN a_6420_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5306 word3.byte3.dff_7.O word3.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5307 VDD a_49620_1704# a_51180_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5308 VDD buf_in30.inv0.O buf_in30.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5309 buf_in18.inv1.O buf_in18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5310 VSS word2.byte3.buf_RE0.O word2.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5311 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5312 a_103080_6578# buf_out16.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5313 a_64560_12850# dec8.and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5314 a_25650_7362# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5315 word4.byte2.dff_4.O word4.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5316 VSS a_22980_6952# a_22940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5317 a_55340_190# a_54550_140# a_55170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5318 a_156900_3442# word3.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5319 a_58380_12184# word8.byte3.cgate0.inv1.O a_57820_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5320 a_155140_10498# a_153300_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5321 a_61650_5912# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5322 buf_sel4.inv1.O buf_sel4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5323 a_62540_11114# word8.byte3.cgate0.inv1.O a_62370_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5324 a_58050_10498# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5325 a_104310_2776# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5326 word3.byte2.tinv7.O word3.byte2.tinv3.EN a_113880_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5327 a_103080_3442# buf_out16.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5328 word2.byte2.dff_4.O word2.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5329 a_25650_4226# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5330 buf_sel5.inv0.O buf_sel5.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5331 a_92280_10500# word7.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5332 VSS a_22980_3816# a_22940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5333 a_14620_11064# a_14950_11904# a_14850_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5334 a_148220_9048# a_147430_8768# a_148050_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5335 VSS buf_in15.inv0.O buf_in15.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5336 VSS word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5337 a_25980_7978# a_25750_8768# a_25420_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5338 VDD a_143500_7928# a_142500_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5339 VDD a_154300_11064# a_153300_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5340 VDD a_121080_6578# a_122640_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5341 a_107910_6462# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5342 a_161730_9598# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5343 a_46020_6578# word5.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5344 word1.byte4.tinv7.O buf_out25.inv0.I a_28020_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5345 VDD a_64020_306# a_65580_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5346 VDD word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5347 a_104920_5912# a_103080_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5348 a_122640_10498# a_122410_9548# a_122080_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5349 VDD a_121080_3442# a_122640_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5350 a_33420_3442# word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5351 a_61750_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5352 VDD word7.byte1.buf_RE1.I word7.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5353 a_107910_3326# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5354 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5355 a_8260_11114# a_6420_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5356 word1.byte1.cgate0.nand0.A word1.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5357 VDD word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5358 VSS word8.byte4.tinv4.I a_17220_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5359 VSS a_126840_680# word1.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5360 a_121080_1704# word2.byte2.tinv5.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5361 VSS a_44580_11764# a_44540_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5362 a_143730_1090# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5363 VSS word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5364 buf_in2.inv1.O buf_in2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5365 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5366 VSS word4.byte2.tinv5.I a_121080_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5367 buf_in24.inv1.O buf_in24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5368 word8.byte3.tinv7.O word8.byte3.tinv0.EN a_42420_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5369 a_122310_10498# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5370 a_101430_190# a_100810_140# a_101320_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5371 word2.gt_re3.I word2.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5372 a_1340_12184# a_550_11904# a_1170_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5373 a_65580_7362# a_65350_6412# a_65020_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5374 a_150700_4792# a_151030_5632# a_150930_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5375 dec8.and4_7.nand0.OUT A0 a_76620_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5376 VDD buf_we2.inv1.O word7.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5377 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5378 VSS a_49620_11112# a_51180_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5379 a_119600_7978# word6.byte2.dff_7.CLK a_119430_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5380 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5381 VSS a_105240_2356# word2.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5382 a_75720_12068# word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5383 VDD a_104080_9548# a_103080_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5384 a_2820_7976# word6.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5385 a_65580_4226# a_65350_3276# a_65020_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5386 VSS a_139900_6412# a_139800_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5387 a_62260_9598# a_60420_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5388 VSS a_122080_4792# a_121080_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5389 a_122640_190# word1.byte2.dff_7.CLK a_122080_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5390 word8.byte3.tinv7.O buf_out20.inv0.I a_56820_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5391 a_73020_9714# word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5392 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5393 a_18550_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5394 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5395 a_57820_4792# word4.byte3.cgate0.inv1.O a_58050_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5396 VSS a_139900_3276# a_139800_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5397 a_103080_4840# word4.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5398 word4.byte2.cgate0.inv1.I word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5399 word8.byte4.dff_2.O word8.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5400 buf_sel6.inv0.O buf_sel6.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5401 VSS a_108840_6952# word5.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5402 a_141020_6462# a_140230_6412# a_140850_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5403 VDD buf_out15.inv0.O buf_out15.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5404 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5405 VSS word3.byte4.tinv6.I a_24420_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5406 VSS a_162660_10088# word7.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5407 VDD word6.byte3.inv_and.O a_75720_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5408 a_101320_7362# a_100380_6462# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5409 word1.byte3.tinv7.O buf_out19.inv0.I a_60420_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5410 a_62580_10088# a_62370_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5411 a_57820_1656# word2.byte3.cgate0.inv1.O a_58050_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5412 a_8580_11764# a_8370_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5413 a_103080_1704# word2.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5414 word2.byte2.cgate0.inv1.I word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5415 VSS buf_out6.inv0.O Do5_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5416 VSS word5.byte3.nand.OUT word5.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5417 a_44260_1090# a_42420_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5418 a_141020_3326# a_140230_3276# a_140850_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5419 VSS a_108840_3816# word3.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5420 a_1170_11114# a_550_11904# a_1060_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5421 a_165430_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5422 a_155460_5492# a_155250_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5423 a_101320_4226# a_100380_3326# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5424 VDD buf_re.inv0.O buf_re.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5425 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5426 a_54550_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5427 a_19340_11114# word8.byte4.cgate0.inv1.O a_19170_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5428 VDD word8.byte2.nand.OUT word8.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5429 VDD a_120_6462# a_780_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5430 buf_in26.inv1.O buf_in26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5431 buf_in8.inv1.O buf_in8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5432 a_155460_2356# a_155250_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5433 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5434 VDD a_144660_680# word1.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5435 a_153300_1704# word2.byte1.tinv3.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5436 a_54550_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5437 a_44580_680# a_44370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5438 Do20_buf buf_out21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5439 buf_in1.inv1.O buf_in1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5440 VSS a_58980_11764# word8.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5441 VDD a_120_3326# a_780_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5442 VSS a_40980_5492# word4.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5443 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5444 buf_sel4.inv1.O buf_sel4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5445 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5446 VSS word6.byte4.nand.OUT word6.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5447 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5448 a_18550_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5449 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5450 VSS word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5451 VSS a_124680_9714# a_126240_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5452 VSS a_58980_8628# word6.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5453 VSS a_20820_6578# a_22380_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5454 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5455 VSS word5.byte2.tinv1.I a_106680_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5456 a_42420_4840# word4.byte3.tinv0.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5457 word5.buf_sel0.O buf_sel5.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X5458 VSS buf_ck.inv0.O CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5459 VSS a_22980_680# word1.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5460 a_140740_190# a_139800_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5461 a_56820_306# word1.byte3.tinv4.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5462 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5463 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5464 a_147940_11114# a_146100_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5465 VDD word5.byte3.tinv1.I a_46020_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5466 word1.byte4.nand.OUT word1.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5467 word2.byte4.dff_4.O word2.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5468 VSS a_20820_3442# a_22380_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5469 a_161500_6412# a_161830_6412# a_161730_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5470 word3.buf_sel0.O buf_sel3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X5471 VDD buf_in11.inv0.O buf_in11.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5472 a_26260_12184# a_24420_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5473 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5474 a_60420_11112# buf_out19.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5475 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5476 VDD word3.byte3.tinv1.I a_46020_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5477 VSS buf_in9.inv0.I buf_in9.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5478 VSS a_61420_9548# a_60420_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5479 word7.byte1.dff_0.O word7.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5480 a_36120_7976# word6.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5481 VDD a_106680_306# a_108240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5482 a_161500_3276# a_161830_3276# a_161730_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5483 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5484 buf_out14.inv1.O buf_out14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5485 word4.byte4.tinv7.O buf_out26.inv0.I a_24420_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5486 buf_in28.inv0.O Di27 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5487 VSS word6.byte1.buf_RE1.I word6.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5488 VDD a_12180_11764# a_12140_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5489 a_50620_9548# a_50950_9548# a_50850_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5490 word7.byte4.tinv7.O buf_out31.inv0.I a_6420_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5491 buf_in17.inv1.O buf_in17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5492 Do4_buf buf_out5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5493 a_144340_2776# a_142500_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5494 VDD a_100480_6412# a_100380_6462# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5495 VSS a_44580_2356# a_44540_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5496 word2.byte4.tinv7.O buf_out26.inv0.I a_24420_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5497 VDD Di19 buf_in20.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5498 a_62540_10498# word7.byte3.cgate0.inv1.O a_62370_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5499 VSS a_15780_8628# a_15740_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5500 VDD a_43420_140# a_42420_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5501 VSS a_116040_6952# a_116000_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5502 VDD a_100480_3276# a_100380_3326# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5503 a_155420_5912# a_154630_5632# a_155250_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5504 a_154530_4842# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5505 a_147940_6462# a_146100_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5506 a_154860_12184# word8.byte1.dff_7.CLK a_154300_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5507 VSS word2.byte3.tinv6.I a_64020_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5508 a_134580_9714# word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5509 a_108240_7362# a_108010_6412# a_107680_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5510 a_33420_5796# word4.byte4.cgate0.nand0.A word4.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5511 word5.byte3.nand.OUT word5.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5512 a_100480_7928# word6.byte2.dff_7.CLK a_100710_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5513 VDD word1.byte1.tinv6.I a_164100_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5514 VSS a_116040_3816# a_116000_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5515 a_112230_4842# a_111610_5632# a_112120_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5516 a_154530_1706# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5517 a_147940_3326# a_146100_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5518 word8.byte4.dff_7.O word8.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5519 VSS word7.gt_re1.O word7.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5520 a_165940_190# a_164100_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5521 a_108240_4226# a_108010_3276# a_107680_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5522 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5523 a_119040_2776# word2.byte2.dff_7.CLK a_118480_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5524 VSS word3.buf_sel0.O word3.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5525 word3.byte3.nand.OUT word3.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5526 a_112230_1706# a_111610_2496# a_112120_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5527 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5528 a_140850_11114# a_140230_11904# a_140740_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5529 a_149700_7976# word6.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5530 a_8260_10498# a_6420_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5531 a_43650_7978# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5532 a_53220_9714# word7.byte3.tinv3.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5533 word6.byte2.tinv7.O buf_out15.inv0.I a_106680_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5534 VDD word6.byte2.buf_RE1.I word6.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5535 VDD a_151860_8628# a_151820_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5536 a_107680_140# a_108010_140# a_107910_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5537 a_140460_6462# word5.byte1.dff_7.CLK a_139900_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5538 word6.byte4.dff_5.O word6.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5539 a_28020_6578# word5.byte4.tinv7.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5540 a_40770_6462# word5.byte3.cgate0.inv1.O a_40660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5541 word5.byte3.dff_3.O word5.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5542 buf_in10.inv1.O buf_in10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5543 a_113880_11112# word8.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5544 a_166260_11764# a_166050_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5545 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5546 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5547 a_140460_3326# word3.byte1.dff_7.CLK a_139900_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5548 a_40770_3326# word3.byte3.cgate0.inv1.O a_40660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5549 word5.byte1.dff_6.O word5.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5550 a_220_7928# word6.byte4.cgate0.inv1.O a_450_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5551 word6.byte1.tinv7.O word6.byte1.tinv3.EN a_153300_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5552 a_43980_190# word1.byte3.cgate0.inv1.O a_43420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5553 word1.byte4.dff_0.O word1.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5554 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5555 buf_in1.inv1.O buf_in1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5556 VSS a_166260_11764# a_166220_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5557 word7.byte4.nand.OUT word7.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5558 buf_in23.inv1.O buf_in23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5559 word3.byte3.dff_3.O word3.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5560 a_55060_4842# a_53220_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5561 VSS word2.byte2.cgate0.inv1.I word2.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5562 VDD a_26580_11764# word8.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5563 word3.byte1.dff_6.O word3.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5564 VDD Di26 buf_in27.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5565 buf_in4.inv1.O buf_in4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5566 a_126630_190# a_126010_140# a_126520_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5567 a_22150_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5568 a_55060_1706# a_53220_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5569 a_17220_11112# buf_out28.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5570 VDD a_155460_5492# word4.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5571 word4.byte2.dff_0.O word4.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5572 VDD A2 dec8.and4_3.nand1.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5573 a_162620_2776# a_161830_2496# a_162450_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5574 buf_sel3.inv1.O buf_sel3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5575 word7.byte4.dff_2.O word7.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5576 a_25750_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5577 VSS a_43420_1656# a_42420_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5578 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5579 a_24420_1704# word2.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5580 VDD a_155460_2356# word2.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5581 word2.byte2.dff_0.O word2.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5582 word8.byte1.tinv7.O buf_out5.inv0.I a_153300_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5583 a_11580_1090# a_11350_140# a_11020_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5584 VSS buf_sel7.inv0.O buf_sel7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5585 a_25750_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5586 a_128280_4840# word4.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5587 a_22940_4842# word4.byte4.cgate0.inv1.O a_22770_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5588 VDD word5.buf_ck1.I word5.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5589 word5.byte2.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5590 VSS word3.byte3.tinv2.I a_49620_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5591 VDD buf_in14.inv0.O buf_in14.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5592 a_1170_9598# a_550_9548# a_1060_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5593 a_126520_7362# a_124680_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5594 a_122640_9048# word6.byte2.dff_7.CLK a_122080_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5595 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5596 word4.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5597 word4.byte3.inv_and.O word4.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5598 a_19340_10498# word7.byte4.cgate0.inv1.O a_19170_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5599 word7.byte4.tinv7.O word7.byte4.tinv3.EN a_13620_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5600 a_128280_1704# word2.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5601 a_22940_1706# word2.byte4.cgate0.inv1.O a_22770_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5602 a_60420_6578# word5.byte3.tinv5.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5603 VDD word3.buf_ck1.I word3.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5604 VDD word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5605 a_126520_4226# a_124680_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5606 a_123200_9598# a_122410_9548# a_123030_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5607 word2.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5608 word2.byte3.inv_and.O word2.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5609 buf_in16.inv1.O buf_in16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5610 VSS a_104080_9548# a_103080_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5611 VDD word6.byte4.tinv4.I a_17220_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5612 a_1380_2356# a_1170_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5613 buf_in7.inv1.O buf_in7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5614 VDD word7.byte4.tinv2.I a_10020_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5615 VDD a_117480_4840# a_119040_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5616 Do19_buf buf_out20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5617 Do0_buf buf_out1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5618 VDD a_19380_8628# a_19340_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5619 VSS a_42420_1704# a_43980_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5620 a_64020_7976# word6.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5621 VDD a_117480_1704# a_119040_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5622 a_106680_4840# word4.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5623 VSS word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5624 word7.byte3.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5625 a_19170_6462# a_18550_6412# a_19060_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5626 a_105200_1090# word1.byte2.dff_7.CLK a_105030_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5627 VSS buf_in22.inv0.O buf_in22.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5628 a_2820_306# word1.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5629 VSS a_13620_7976# a_15180_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5630 a_20820_7976# word6.byte4.tinv5.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5631 a_108520_11114# a_106680_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5632 a_147940_10498# a_146100_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5633 a_158850_7978# a_158230_8768# a_158740_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5634 word5.byte2.tinv7.O buf_out11.inv0.I a_121080_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5635 a_55170_4842# word4.byte3.cgate0.inv1.O a_55060_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5636 buf_sel1.inv0.I dec8.and4_0.nand1.OUT a_65100_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5637 VSS a_46020_6578# a_47580_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5638 VDD word4.byte4.tinv1.I a_6420_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5639 VDD a_22980_8628# word6.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5640 a_67620_5796# word4.byte3.tinv7.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5641 a_19170_3326# a_18550_3276# a_19060_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5642 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5643 word4.byte3.dff_7.O word4.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5644 VDD a_156900_6578# a_158460_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5645 a_154300_7928# a_154630_8768# a_154530_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5646 a_115830_190# word1.byte2.dff_7.CLK a_115720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5647 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.latch0.I0.O a_131700_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5648 word3.byte2.tinv7.O buf_out11.inv0.I a_121080_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5649 VDD word2.byte4.tinv1.I a_6420_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5650 VSS a_46020_3442# a_47580_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5651 a_43420_4792# word4.byte3.cgate0.inv1.O a_43650_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5652 VDD word5.gt_re1.O word5.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5653 VDD word1.byte3.inv_and.O a_75720_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5654 VDD word4.buf_ck1.I word4.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5655 word6.byte1.inv_and.O word6.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5656 VDD a_8580_5492# a_8540_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5657 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5658 VDD a_156900_3442# a_158460_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5659 word3.gt_re0.OUT buf_sel3.inv1.O a_82020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5660 a_43650_12184# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5661 a_61980_11114# a_61750_11904# a_61420_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5662 a_108800_12184# a_108010_11904# a_108630_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5663 a_151030_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5664 VDD a_12180_10088# a_12140_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5665 a_43420_1656# word2.byte3.cgate0.inv1.O a_43650_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5666 word7.byte1.dff_7.O word7.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5667 a_105240_6952# a_105030_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5668 VDD word2.buf_ck1.I word2.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5669 VDD word3.gt_re1.O word3.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5670 VDD a_8580_2356# a_8540_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5671 a_49620_4840# buf_out22.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5672 VDD a_149700_7976# a_151260_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5673 a_158130_190# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5674 VDD buf_in27.inv0.O buf_in27.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5675 word5.byte4.tinv7.O word5.byte4.tinv5.EN a_20820_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5676 VSS a_22980_5492# a_22940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5677 a_43420_11064# word8.byte3.cgate0.inv1.O a_43650_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5678 a_105240_3816# a_105030_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5679 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5680 a_156900_9714# buf_out4.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5681 a_49620_1704# buf_out22.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5682 Do24_buf buf_out25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5683 VDD a_125680_6412# a_124680_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5684 VDD a_62580_6952# word5.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5685 a_14850_9598# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5686 a_780_9048# word6.byte4.cgate0.inv1.O a_220_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5687 a_1170_4842# a_550_5632# a_1060_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5688 VSS word8.byte4.cgate0.nand0.A a_35760_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5689 word1.byte1.dff_2.O word1.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5690 VSS word2.byte1.buf_RE1.I word2.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5691 word6.gt_re3.I word6.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5692 a_6420_306# word1.byte4.tinv1.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5693 VDD a_125680_3276# a_124680_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5694 a_107910_5912# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5695 a_125680_140# word1.byte2.dff_7.CLK a_125910_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5696 a_7980_2776# word2.byte4.cgate0.inv1.O a_7420_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5697 VDD a_62580_3816# word3.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5698 VSS buf_out19.inv0.O Do18_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5699 a_149700_306# word1.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5700 a_1170_1706# a_550_2496# a_1060_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5701 word2.byte1.nand.B word2.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5702 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5703 a_101430_11114# a_100810_11904# a_101320_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5704 a_140850_9598# a_140230_9548# a_140740_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5705 VSS a_110280_9714# a_111840_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5706 a_117480_9714# word7.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5707 word8.byte1.dff_2.O word8.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5708 VDD word7.buf_ck1.I word7.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5709 a_162060_2776# word2.byte1.dff_7.CLK a_161500_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5710 word8.byte4.cgate0.inv1.I word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5711 a_26260_6462# a_24420_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5712 a_62370_1706# word2.byte3.cgate0.inv1.O a_62260_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5713 a_129540_9714# word7.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5714 word4.byte4.tinv7.O word4.byte4.tinv7.EN a_28020_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5715 a_4050_6462# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5716 VSS word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5717 VSS word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5718 a_122410_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5719 a_126840_11764# a_126630_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5720 a_166260_10088# a_166050_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5721 a_126240_7978# a_126010_8768# a_125680_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5722 a_36120_1092# word1.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5723 a_22380_4842# a_22150_5632# a_21820_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5724 a_26260_3326# a_24420_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5725 a_4050_3326# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5726 a_165660_6462# word5.byte1.dff_7.CLK a_165100_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5727 buf_in16.inv1.O buf_in16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5728 word6.byte3.dff_1.O word6.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5729 a_65970_6462# word5.byte3.cgate0.inv1.O a_65860_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5730 VSS a_101640_11764# a_101600_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5731 a_42420_3442# word3.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5732 buf_in9.inv1.O buf_in9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5733 a_26580_6952# a_26370_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5734 VDD word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5735 word8.byte1.dff_5.O word8.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5736 a_22380_1706# a_22150_2496# a_21820_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5737 VDD a_26580_10088# word7.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5738 VSS word8.byte2.buf_RE1.I word8.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5739 a_165660_3326# word3.byte1.dff_7.CLK a_165100_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5740 word4.byte4.tinv7.O buf_out30.inv0.I a_10020_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5741 a_65970_3326# word3.byte3.cgate0.inv1.O a_65860_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5742 VSS word6.byte2.tinv6.I a_124680_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5743 a_26580_3816# a_26370_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5744 VSS a_139900_4792# a_139800_4842# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5745 a_11970_190# word1.byte4.cgate0.inv1.O a_11860_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5746 buf_in3.inv1.O buf_in3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5747 a_54780_9598# word7.byte3.cgate0.inv1.O a_54220_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5748 a_66140_6462# a_65350_6412# a_65970_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5749 a_148260_2356# a_148050_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5750 word2.byte4.tinv7.O buf_out30.inv0.I a_10020_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5751 VDD buf_out30.inv0.O Do29_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5752 buf_in26.inv1.O buf_in26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5753 buf_in3.inv1.O buf_in3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5754 a_39180_12068# buf_we1.inv1.O word8.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5755 a_104310_7362# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5756 a_47350_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5757 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5758 a_118810_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5759 VSS a_101640_6952# a_101600_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5760 a_67620_10500# word7.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5761 word4.byte2.dff_7.O word4.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5762 a_141020_5912# a_140230_5632# a_140850_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5763 VSS a_108840_5492# word4.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5764 a_18780_11114# a_18550_11904# a_18220_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5765 word8.byte2.tinv7.O buf_out13.inv0.I a_113880_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5766 VSS a_125680_7928# a_124680_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5767 a_66140_3326# a_65350_3276# a_65970_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5768 a_18550_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5769 a_104310_4226# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5770 buf_in32.inv1.O buf_in32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5771 VDD buf_in18.inv0.O buf_in18.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5772 a_49620_1704# word2.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5773 VSS a_101640_3816# a_101600_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5774 word2.byte2.dff_7.O word2.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5775 a_149700_306# word1.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5776 a_159020_9048# a_158230_8768# a_158850_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5777 a_157900_7928# word6.byte1.dff_7.CLK a_158130_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5778 VSS buf_sel8.inv0.O buf_sel8.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5779 VSS word7.byte3.buf_RE0.O word7.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5780 a_82020_9714# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5781 a_124680_6578# word5.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5782 word4.byte3.tinv7.O word4.byte3.tinv5.EN a_60420_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5783 a_108840_10088# a_108630_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5784 VDD word1.byte2.buf_RE1.I word1.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5785 word1.byte2.tinv7.O buf_out15.inv0.I a_106680_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5786 a_11250_11114# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5787 VSS word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5788 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5789 VSS word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5790 word5.byte3.cgate0.nand0.A word5.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5791 a_47350_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5792 VDD a_6420_4840# a_7980_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5793 buf_in15.inv1.O buf_in15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5794 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5795 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5796 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5797 a_11020_1656# a_11350_2496# a_11250_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5798 word4.byte3.cgate0.inv1.I word4.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5799 a_154630_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5800 VSS a_25420_6412# a_24420_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5801 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5802 buf_out9.inv1.O buf_out9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5803 VSS a_66180_10088# word7.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5804 VDD a_6420_1704# a_7980_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5805 word2.byte3.cgate0.inv1.I word2.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5806 a_19060_190# a_17220_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5807 a_40660_4842# a_39720_4842# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5808 VSS a_20820_4840# a_22380_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5809 a_14620_6412# a_14950_6412# a_14850_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5810 VSS a_25420_3276# a_24420_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5811 a_55060_11114# a_53220_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5812 VSS word6.byte1.tinv4.I a_156900_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5813 a_108520_10498# a_106680_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5814 VDD a_105240_6952# word5.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5815 word6.byte4.cgate0.nand0.A word6.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5816 a_40660_1706# a_39720_1706# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5817 a_14620_3276# a_14950_3276# a_14850_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5818 a_161500_4792# a_161830_5632# a_161730_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5819 VDD a_10020_11112# a_11580_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5820 a_46020_7976# word6.byte3.tinv1.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5821 a_151860_8628# a_151650_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5822 VDD a_141060_5492# word4.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5823 VDD a_48180_680# word1.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5824 a_40980_5492# a_40770_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5825 VDD buf_in2.inv0.O buf_in2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5826 VDD a_105240_3816# word3.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5827 a_146100_6578# buf_out7.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5828 dec8.and4_2.nand0.OUT dec8.and4_6.nand0.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5829 VSS word5.byte4.dff_0.O_bar a_2820_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5830 VSS a_116040_2356# word2.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5831 VSS word4.byte1.nand.B a_39180_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5832 VDD a_141060_2356# word2.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X5833 a_61980_10498# a_61750_9548# a_61420_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5834 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5835 a_147330_2776# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5836 a_24420_11112# word8.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5837 a_40980_2356# a_40770_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5838 a_151030_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5839 word3.byte1.tinv7.O word3.byte1.tinv4.EN a_156900_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5840 a_146100_3442# buf_out7.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5841 a_62540_190# a_61750_140# a_62370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5842 VSS word3.byte2.tinv0.I a_103080_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5843 a_113880_4840# word4.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5844 VDD buf_sel6.inv0.O buf_sel6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5845 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5846 a_158850_11114# a_158230_11904# a_158740_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5847 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5848 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5849 a_11970_11114# word8.byte4.cgate0.inv1.O a_11860_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5850 a_165330_12184# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5851 a_43420_9548# word7.byte3.cgate0.inv1.O a_43650_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5852 VDD word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5853 word6.byte3.dff_2.O word6.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5854 word1.byte2.tinv7.O word1.byte2.tinv4.EN a_117480_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5855 word5.byte1.nand.B word5.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5856 a_113880_1704# word2.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5857 a_117480_9714# buf_out12.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5858 VDD word1.byte4.tinv4.I a_17220_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5859 VSS a_116040_5492# a_116000_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5860 a_108630_6462# word5.byte2.dff_7.CLK a_108520_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5861 word8.byte3.dff_4.O word8.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5862 a_147940_5912# a_146100_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5863 a_162450_9598# word7.byte1.dff_7.CLK a_162340_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5864 word5.byte3.tinv7.O word5.byte3.tinv1.EN a_46020_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5865 a_165100_11064# word8.byte1.dff_7.CLK a_165330_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5866 VDD buf_in32.inv0.O buf_in32.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5867 Do7_buf buf_out8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5868 a_108630_3326# word3.byte2.dff_7.CLK a_108520_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5869 VDD a_103080_4840# a_104640_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5870 a_164100_1704# word2.byte1.tinv6.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5871 a_40050_9598# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X5872 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5873 VDD a_43420_9548# a_42420_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5874 a_123240_8628# a_123030_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5875 a_55380_680# a_55170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5876 VDD Di28 buf_in29.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5877 word8.byte1.tinv7.O word8.byte1.tinv4.EN a_156900_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5878 VSS a_65020_140# a_64020_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5879 buf_re.inv1.O buf_re.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5880 VSS word8.byte4.buf_RE0.O word8.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5881 a_101430_9598# a_100810_9548# a_101320_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5882 VDD a_103080_1704# a_104640_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5883 a_2820_9714# buf_out32.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X5884 VSS buf_in18.inv0.O buf_in18.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5885 VSS word4.byte1.tinv6.I a_164100_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5886 a_144450_190# a_143830_140# a_144340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5887 word2.byte3.cgate0.inv1.O word2.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5888 VSS a_164100_11112# a_165660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5889 a_140460_5912# word4.byte1.dff_7.CLK a_139900_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5890 CLK buf_ck.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5891 word5.byte4.dff_4.O word5.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5892 a_40770_4842# word4.byte3.cgate0.inv1.O a_40660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5893 a_19060_9048# a_17220_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5894 VSS word2.byte4.buf_RE0.O word2.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5895 VDD word7.gt_re1.O word7.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5896 a_126840_10088# a_126630_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X5897 word4.byte3.dff_3.O word4.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5898 VSS buf_sel4.inv0.O buf_sel4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5899 VSS a_148260_2356# word2.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5900 word1.byte1.inv_and.O word1.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5901 VSS a_119640_8628# word6.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X5902 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5903 word3.byte4.dff_4.O word3.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5904 VDD word5.byte3.tinv4.I a_56820_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5905 a_158460_9048# word6.byte1.dff_7.CLK a_157900_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5906 word7.byte1.dff_5.O word7.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5907 word6.byte4.tinv7.O buf_out32.inv0.I a_2820_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5908 a_58770_7978# word6.byte3.cgate0.inv1.O a_58660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5909 VDD a_165100_4792# a_164100_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5910 a_47580_4842# a_47350_5632# a_47020_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5911 a_146100_4840# word4.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5912 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5913 a_67620_3442# word3.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5914 VDD word3.byte3.tinv4.I a_56820_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5915 word7.byte1.dff_3.O word7.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5916 a_25750_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5917 a_15740_2776# a_14950_2496# a_15570_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5918 a_144340_7362# a_142500_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5919 VDD a_44580_6952# a_44540_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5920 VDD a_165100_1656# a_164100_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5921 a_47580_1706# a_47350_2496# a_47020_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5922 a_146100_1704# word2.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5923 a_24420_3442# word3.byte4.tinv6.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5924 buf_in11.inv1.O buf_in11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5925 VDD word4.byte4.cgate0.nand0.A a_35760_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5926 VDD word6.byte1.cgate0.nand0.B word6.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5927 VSS a_123240_2356# a_123200_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5928 VDD word8.byte1.cgate0.nand0.B word8.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5929 a_144340_4226# a_142500_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5930 a_25750_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X5931 buf_in11.inv0.O buf_in11.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X5932 a_18780_10498# a_18550_9548# a_18220_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5933 VDD word7.byte4.tinv7.I a_28020_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5934 VDD a_54220_7928# a_53220_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X5935 VDD a_44580_3816# a_44540_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5936 buf_in25.inv1.O buf_in25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5937 VSS a_3820_140# a_2820_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5938 VDD word2.byte4.cgate0.nand0.A a_35760_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5939 buf_in7.inv1.O buf_in7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5940 VSS a_126840_6952# a_126800_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5941 VSS buf_in24.inv0.O buf_in24.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5942 a_111280_140# word1.byte2.dff_7.CLK a_111510_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X5943 VSS buf_in17.inv0.O buf_in17.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5944 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5945 a_119040_7362# a_118810_6412# a_118480_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5946 VSS word1.byte4.tinv7.I a_28020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5947 VSS a_143500_4792# a_142500_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X5948 buf_in31.inv1.O buf_in31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5949 a_160500_11112# word8.byte1.tinv5.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5950 a_123030_4842# a_122410_5632# a_122920_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5951 VSS a_126840_3816# a_126800_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5952 a_11250_10498# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5953 VSS word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5954 a_11860_6462# a_10020_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5955 a_54450_1090# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5956 a_119040_4226# a_118810_3276# a_118480_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5957 a_47350_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5958 a_115720_9598# a_113880_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5959 a_122310_7978# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X5960 a_123030_1706# a_122410_2496# a_122920_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5961 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5962 VSS word5.byte1.tinv2.I a_149700_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5963 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5964 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5965 buf_sel2.inv0.O buf_sel2.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5966 VDD a_162660_680# a_162620_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5967 a_64020_9714# word7.byte3.tinv6.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5968 a_111840_7978# a_111610_8768# a_111280_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5969 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5970 a_106680_6578# word5.byte2.tinv1.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5971 a_11860_3326# a_10020_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5972 a_143830_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5973 VDD word5.buf_sel0.O word5.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5974 VDD word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5975 a_64020_306# word1.byte3.tinv6.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X5976 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5977 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5978 buf_out15.inv1.O buf_out15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5979 a_7420_9548# a_7750_9548# a_7650_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5980 VDD word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5981 a_12180_6952# a_11970_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5982 VSS buf_in32.inv0.O buf_in32.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5983 a_55060_10498# a_53220_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5984 VSS word5.byte3.buf_RE0.O word5.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5985 VDD word3.buf_sel0.O word3.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5986 VDD word8.byte3.cgate0.nand0.A word8.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X5987 a_22150_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X5988 a_107680_6412# a_108010_6412# a_107910_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X5989 VDD word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X5990 a_12180_3816# a_11970_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X5991 buf_re.inv1.O buf_re.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X5992 word6.byte4.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X5993 a_65860_4842# a_64020_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X5994 VSS a_46020_4840# a_47580_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X5995 a_101040_12184# word8.byte2.dff_7.CLK a_100480_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5996 VDD a_10020_9714# a_11580_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X5997 a_51740_6462# a_50950_6412# a_51570_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5998 a_126240_12184# word8.byte2.dff_7.CLK a_125680_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X5999 VSS a_4980_2356# word2.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6000 Do3_buf buf_out4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6001 a_107680_3276# a_108010_3276# a_107910_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6002 a_22150_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6003 a_2820_4840# word4.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6004 a_162620_7362# word5.byte1.dff_7.CLK a_162450_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6005 a_1340_1090# word1.byte4.cgate0.inv1.O a_1170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6006 a_65860_1706# a_64020_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6007 VSS buf_in1.inv0.O buf_in1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6008 a_51740_3326# a_50950_3276# a_51570_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6009 VSS a_146100_9714# a_147660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6010 a_104410_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6011 word1.byte4.tinv7.O word1.byte4.tinv6.EN a_24420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6012 a_103080_1704# word2.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6013 a_95160_2660# word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6014 a_66180_5492# a_65970_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6015 VSS a_159060_6952# a_159020_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6016 a_162620_4226# word3.byte1.dff_7.CLK a_162450_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6017 VDD buf_out19.inv0.I buf_out19.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X6018 a_119430_11114# a_118810_11904# a_119320_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6019 a_158850_9598# a_158230_9548# a_158740_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6020 VSS word6.byte4.buf_RE0.O word6.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6021 a_100710_12184# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6022 VDD word7.byte1.cgate0.nand0.B word7.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6023 VSS word4.byte3.inv_and.O a_75720_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6024 dec8.and4_4.nand1.OUT A2 a_71760_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6025 a_155250_4842# a_154630_5632# a_155140_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6026 a_101600_4842# word4.byte2.dff_7.CLK a_101430_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6027 a_146100_11112# word8.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6028 a_143500_7928# word6.byte1.dff_7.CLK a_143730_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6029 a_66180_2356# a_65970_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6030 VSS a_159060_3816# a_159020_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6031 a_104410_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6032 VDD a_123240_8628# word6.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6033 VDD a_19380_5492# word4.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6034 a_134580_9714# word7.byte1.cgate0.nand0.A word7.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6035 VSS word3.byte2.tinv7.I a_128280_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6036 VDD CLK word5.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6037 dec8.and4_3.nand1.A A2 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6038 VSS word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6039 VDD buf_sel3.inv0.O buf_sel3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6040 word7.byte3.dff_4.O word7.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6041 word5.byte4.dff_2.O word5.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6042 a_101600_1706# word2.byte2.dff_7.CLK a_101430_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6043 a_100480_11064# word8.byte2.dff_7.CLK a_100710_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6044 VSS a_48180_10088# a_48140_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6045 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6046 a_155250_1706# a_154630_2496# a_155140_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6047 a_1380_6952# a_1170_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6048 VDD a_19380_2356# word2.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6049 a_125680_11064# word8.byte2.dff_7.CLK a_125910_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6050 a_165100_9548# word7.byte1.dff_7.CLK a_165330_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6051 a_149700_7976# buf_out6.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6052 a_140230_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6053 buf_in11.inv1.O buf_in11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6054 VSS a_119640_11764# a_119600_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6055 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6056 VDD CLK word3.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6057 word8.byte1.dff_3.O word8.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6058 word3.byte4.dff_2.O word3.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6059 buf_in16.inv1.O buf_in16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6060 VSS a_114880_9548# a_113880_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6061 a_1380_3816# a_1170_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6062 word8.byte2.tinv7.O word8.byte2.tinv4.EN a_117480_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6063 VSS a_51780_10088# word7.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6064 a_15180_2776# word2.byte4.cgate0.inv1.O a_14620_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6065 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6066 a_151860_11764# a_151650_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6067 VDD a_42420_6578# a_43980_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6068 a_39820_7928# a_40150_8768# a_40050_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6069 word1.byte2.nand.OUT buf_we3.inv1.O a_90120_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6070 a_114880_140# a_115210_140# a_115110_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6071 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6072 VSS Di27 buf_in28.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6073 VSS buf_out14.inv0.O buf_out14.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6074 VSS word6.byte1.tinv0.I a_142500_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6075 VDD a_165100_9548# a_164100_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6076 VDD a_42420_3442# a_43980_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6077 a_26260_5912# a_24420_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6078 VSS a_12180_11764# word8.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6079 a_18780_6462# word5.byte4.cgate0.inv1.O a_18220_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6080 VSS a_53220_1704# a_54780_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6081 a_4050_5912# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6082 VSS word6.byte2.inv_and.O a_92280_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6083 a_11250_6462# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6084 a_36120_306# word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6085 VSS a_4980_11764# a_4940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6086 a_116000_1090# word1.byte2.dff_7.CLK a_115830_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6087 a_18780_3326# word3.byte4.cgate0.inv1.O a_18220_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6088 a_165660_5912# word4.byte1.dff_7.CLK a_165100_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6089 VDD buf_out3.inv0.O Do2_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6090 word8.byte4.tinv7.O word8.byte4.tinv0.EN a_2820_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6091 word4.byte1.dff_1.O word4.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6092 a_65970_4842# word4.byte3.cgate0.inv1.O a_65860_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6093 a_56820_11112# word8.byte3.tinv4.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6094 a_11250_3326# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6095 a_26580_5492# a_26370_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6096 a_122080_4792# word4.byte2.dff_7.CLK a_122310_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6097 VSS word1.byte1.cgate0.nand0.B a_134580_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6098 VSS word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6099 word2.byte1.dff_1.O word2.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6100 a_36120_5796# word4.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6101 a_22770_7978# a_22150_8768# a_22660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6102 word2.byte4.tinv7.O word2.byte4.tinv6.EN a_24420_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6103 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6104 a_122080_1656# word2.byte2.dff_7.CLK a_122310_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6105 word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.latch0.I0.O a_92280_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6106 a_66140_5912# a_65350_5632# a_65970_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6107 a_142500_6578# word5.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6108 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6109 a_65250_4842# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6110 VDD a_160500_306# a_162060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6111 word3.byte4.inv_and.O word3.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6112 a_92280_6578# word5.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6113 VSS word5.byte2.buf_RE1.I word5.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6114 VSS a_101640_5492# a_101600_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6115 VSS a_126840_11764# word8.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6116 a_65250_1706# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6117 VDD word6.byte3.tinv5.I a_60420_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6118 VSS a_104080_11064# a_103080_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6119 a_124680_9714# word7.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6120 a_166220_9598# a_165430_9548# a_166050_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6121 VSS buf_in10.inv0.O buf_in10.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6122 a_7980_7362# a_7750_6412# a_7420_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6123 a_47860_11114# a_46020_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6124 VSS a_119640_8628# a_119600_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6125 a_140130_190# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6126 a_108520_4842# a_106680_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6127 buf_in27.inv1.O buf_in27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6128 a_17220_7976# buf_out28.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6129 a_162340_7978# a_160500_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6130 VDD a_62580_8628# a_62540_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6131 a_51180_6462# word5.byte3.cgate0.inv1.O a_50620_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6132 word7.byte1.tinv7.O buf_out6.inv0.I a_149700_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6133 a_7980_4226# a_7750_3276# a_7420_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6134 a_4660_9598# a_2820_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6135 buf_in30.inv1.O buf_in30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6136 a_162060_7362# a_161830_6412# a_161500_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6137 a_62370_6462# a_61750_6412# a_62260_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6138 a_108520_1706# a_106680_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6139 a_149700_4840# word4.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6140 VDD a_118480_11064# a_117480_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6141 VDD buf_in21.inv0.O buf_in21.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6142 a_35760_12068# word8.byte1.cgate0.nand0.B word8.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6143 a_148220_1090# word1.byte1.dff_7.CLK a_148050_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6144 a_51180_3326# word3.byte3.cgate0.inv1.O a_50620_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6145 word6.byte3.tinv7.O word6.byte3.tinv6.EN a_64020_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6146 a_40940_12184# a_40150_11904# a_40770_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6147 a_162060_4226# a_161830_3276# a_161500_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6148 word4.byte2.tinv7.O word4.byte2.tinv1.EN a_106680_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6149 VSS word4.byte2.buf_RE1.I word4.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6150 a_66140_12184# a_65350_11904# a_65970_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6151 a_62370_3326# a_61750_3276# a_62260_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6152 word5.byte1.tinv7.O buf_out2.inv0.I a_164100_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6153 VSS buf_sel3.inv0.O buf_sel3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6154 a_104410_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6155 VDD word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6156 word7.byte1.nand.B word7.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6157 a_143830_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6158 VDD word5.byte2.tinv2.I a_110280_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6159 word1.byte4.tinv7.O buf_out32.inv0.I a_2820_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6160 a_131700_306# word1.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6161 a_4980_10088# a_4770_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6162 VSS a_139900_140# a_139800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6163 a_132960_6578# word5.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6164 a_6420_4840# buf_out31.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6165 dec8.and4_3.nand1.OUT dec8.and4_3.nand1.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6166 a_35760_9714# word7.byte1.cgate0.nand0.B word7.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6167 word6.byte2.dff_6.O word6.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6168 word3.byte1.tinv7.O buf_out2.inv0.I a_164100_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6169 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6170 a_14620_4792# a_14950_5632# a_14850_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6171 a_121080_3442# word3.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6172 VDD word3.byte2.tinv2.I a_110280_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6173 VDD a_150700_4792# a_149700_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6174 a_131700_4840# word4.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6175 VDD word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6176 a_123030_190# word1.byte2.dff_7.CLK a_122920_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6177 a_6420_1704# buf_out31.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6178 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B a_132960_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6179 VDD word1.byte1.cgate0.nand0.B word1.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6180 VDD word4.buf_ck1.I word4.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6181 VDD a_150700_1656# a_149700_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6182 a_131700_1704# word2.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6183 a_10020_3442# word3.byte4.tinv2.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6184 a_148260_6952# a_148050_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6185 buf_out12.inv1.O buf_out12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6186 VDD word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6187 a_93540_4840# word4.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6188 a_47350_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6189 word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.latch0.I0.ENB a_75720_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6190 a_44540_9048# a_43750_8768# a_44370_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6191 VSS a_156900_306# a_158460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6192 a_151030_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6193 a_48180_11764# a_47970_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6194 VDD word2.buf_ck1.I word2.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6195 VSS word5.byte4.tinv2.I a_10020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6196 a_20820_7976# word6.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6197 a_126010_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6198 a_148260_3816# a_148050_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6199 a_40770_11114# a_40150_11904# a_40660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6200 a_165330_190# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6201 a_93540_1704# word2.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6202 a_47350_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6203 VDD buf_out10.inv0.O buf_out10.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6204 a_151030_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6205 a_119430_9598# a_118810_9548# a_119320_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6206 a_141060_8628# a_140850_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6207 VSS buf_out1.inv0.O Do0_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6208 a_40150_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6209 word6.byte1.cgate0.inv1.I word6.byte1.cgate0.nand0.A a_134580_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6210 a_128280_2660# word2.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6211 Do29_buf buf_out30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6212 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6213 a_100810_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6214 word2.byte2.nand.OUT buf_we3.inv1.O a_90120_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6215 word2.byte3.inv_and.O word2.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6216 a_108630_4842# word4.byte2.dff_7.CLK a_108520_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6217 a_100480_9548# word7.byte2.dff_7.CLK a_100710_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6218 VSS word7.byte1.tinv5.I a_160500_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6219 a_126800_4842# word4.byte2.dff_7.CLK a_126630_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6220 VSS a_66180_680# word1.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6221 a_156900_306# word1.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6222 a_125680_9548# word7.byte2.dff_7.CLK a_125910_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6223 VDD a_44580_5492# word4.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6224 a_21820_140# a_22150_140# a_22050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6225 VSS word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6226 a_73020_12068# word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6227 a_11020_6412# word5.byte4.cgate0.inv1.O a_11250_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6228 VDD buf_sel4.inv0.O buf_sel4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6229 word8.byte2.dff_3.O word8.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6230 VSS a_3820_9548# a_2820_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6231 word7.byte1.dff_3.O word7.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6232 a_126800_1706# word2.byte2.dff_7.CLK a_126630_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6233 word7.byte2.tinv7.O word7.byte2.tinv4.EN a_117480_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6234 VSS word7.byte1.nand.OUT word7.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6235 VSS word4.byte4.tinv4.I a_17220_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6236 VDD a_44580_2356# word2.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6237 VDD word8.byte4.tinv5.I a_20820_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6238 a_92280_10500# word7.byte2.cgate0.latch0.I0.ENB word7.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6239 a_165430_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6240 buf_sel5.inv1.O buf_sel5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6241 VDD word8.byte3.tinv1.I a_46020_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6242 a_11020_3276# word3.byte4.cgate0.inv1.O a_11250_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6243 buf_in15.inv1.O buf_in15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6244 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6245 a_73020_3442# word3.byte3.cgate0.nand0.A word3.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6246 VDD word4.gt_re1.O word4.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6247 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6248 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6249 VDD word4.byte4.buf_RE0.O word4.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6250 word1.byte4.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6251 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6252 a_65020_7928# a_65350_8768# a_65250_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6253 VDD word2.gt_re1.O word2.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6254 buf_in13.inv0.O buf_in13.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6255 VSS word1.byte2.tinv0.I a_103080_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6256 word3.byte3.tinv7.O word3.byte3.tinv0.EN a_42420_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6257 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6258 buf_in27.inv1.O buf_in27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6259 VDD word6.byte1.cgate0.nand0.B word6.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6260 VSS word6.byte1.tinv7.I a_167700_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6261 VSS a_141060_2356# a_141020_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6262 VDD word2.byte4.buf_RE0.O word2.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6263 VDD a_18220_4792# a_17220_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6264 VSS word2.byte4.tinv1.I a_6420_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6265 VDD a_116040_6952# word5.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6266 a_124680_7976# word6.byte2.tinv6.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6267 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6268 word7.byte3.tinv7.O buf_out23.inv0.I a_46020_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6269 VSS buf_out30.inv0.I buf_out30.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X6270 a_119640_5492# a_119430_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6271 VDD a_58980_680# word1.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6272 VDD a_18220_1656# a_17220_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6273 a_147330_7362# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6274 VDD a_60420_7976# a_61980_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6275 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6276 a_61750_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6277 a_75360_8932# word6.byte1.cgate0.nand0.B word6.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6278 VSS word2.buf_ck1.I word2.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6279 VSS a_144660_6952# a_144620_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6280 VDD buf_in2.inv0.O buf_in2.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6281 VDD a_116040_3816# word3.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6282 word4.byte1.inv_and.O word4.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6283 buf_in24.inv0.O Di23 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6284 VSS a_4980_680# word1.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6285 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6286 VSS a_100380_7978# a_101040_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6287 a_119640_2356# a_119430_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6288 VSS word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6289 a_147330_4226# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6290 VDD CLK word7.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6291 a_140850_4842# a_140230_5632# a_140740_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6292 VSS dec8.and4_7.nand0.OUT buf_sel8.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6293 VSS a_144660_3816# a_144620_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6294 a_47020_140# a_47350_140# a_47250_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6295 a_49620_1704# word2.byte3.tinv2.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6296 a_147660_7978# a_147430_8768# a_147100_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6297 Do16_buf buf_out17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6298 a_47970_7978# a_47350_8768# a_47860_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6299 a_149700_306# buf_out6.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6300 a_115830_1706# word2.byte2.dff_7.CLK a_115720_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6301 a_140130_7978# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6302 a_140850_1706# a_140230_2496# a_140740_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6303 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6304 a_167700_6578# word5.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6305 word6.byte3.dff_5.O word6.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6306 a_148220_190# a_147430_140# a_148050_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6307 word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.latch0.I0.O a_75720_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6308 word7.gt_re1.O word7.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6309 VDD word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6310 VDD word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6311 word5.byte2.tinv7.O word5.byte2.tinv6.EN a_124680_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6312 VSS a_126840_5492# a_126800_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6313 a_47860_10498# a_46020_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6314 buf_sel6.inv1.O buf_sel6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6315 VSS word7.byte4.tinv7.I a_28020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6316 word3.byte4.cgate0.inv1.I word3.byte4.cgate0.nand0.A a_33420_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6317 a_15780_11764# a_15570_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6318 a_48140_7978# word6.byte3.cgate0.inv1.O a_47970_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6319 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6320 VSS word1.byte2.tinv7.I a_128280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6321 a_118710_9598# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6322 VSS word1.byte2.buf_RE1.I word1.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6323 VDD word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6324 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6325 VDD a_65020_11064# a_64020_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6326 a_119040_12184# word8.byte2.dff_7.CLK a_118480_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6327 a_162340_11114# a_160500_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6328 VDD a_15780_680# a_15740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6329 a_11860_5912# a_10020_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6330 Do29_buf buf_out30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6331 VSS buf_in26.inv0.O buf_in26.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6332 a_26260_190# a_24420_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6333 a_58660_2776# a_56820_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6334 a_104410_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6335 VDD a_148260_6952# word5.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6336 VDD buf_in8.inv0.O buf_in8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6337 VDD buf_out21.inv0.I buf_out21.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X6338 VDD buf_in1.inv0.O buf_in1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6339 a_12180_5492# a_11970_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6340 a_118710_12184# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6341 a_162620_12184# a_161830_11904# a_162450_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6342 a_49620_9714# buf_out22.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6343 VDD a_148260_3816# word3.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6344 VSS buf_in32.inv0.O buf_in32.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6345 VSS buf_sel4.inv0.O buf_sel4.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6346 VDD word8.byte1.buf_RE1.I word8.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6347 VSS a_159060_2356# word2.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6348 a_58980_2356# a_58770_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6349 a_107680_4792# a_108010_5632# a_107910_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6350 VSS word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6351 a_64020_11112# word8.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6352 a_15740_7362# word5.byte4.cgate0.inv1.O a_15570_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6353 VDD buf_ck.inv0.O CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6354 VSS word8.buf_sel0.O word8.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6355 a_2820_6578# word5.byte4.tinv0.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6356 word1.byte4.dff_5.O word1.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6357 a_161730_9048# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6358 a_112120_6462# a_110280_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6359 word2.byte4.tinv7.O word2.byte4.tinv2.EN a_10020_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6360 a_144450_11114# word8.byte1.dff_7.CLK a_144340_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6361 VSS word3.byte1.tinv1.I a_146100_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6362 a_156900_4840# word4.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6363 a_118480_11064# word8.byte2.dff_7.CLK a_118710_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6364 a_51740_5912# a_50950_5632# a_51570_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6365 word7.gt_re3.I word7.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6366 a_50850_4842# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6367 a_36120_11112# word8.byte4.cgate0.latch0.I0.ENB word8.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6368 VDD a_123240_6952# a_123200_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6369 VSS word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6370 VSS a_12180_2356# word2.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6371 a_15740_4226# word3.byte4.cgate0.inv1.O a_15570_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6372 a_11350_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6373 word4.byte2.tinv7.O buf_out13.inv0.I a_113880_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6374 a_112120_3326# a_110280_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6375 VSS word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6376 VDD word1.byte3.tinv5.I a_60420_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6377 a_156900_1704# word2.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6378 a_40770_9598# a_40150_9548# a_40660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6379 buf_in11.inv1.O buf_in11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6380 a_4050_12184# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6381 a_3820_6412# a_4150_6412# a_4050_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6382 a_18450_190# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6383 a_50850_1706# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6384 VDD a_123240_3816# a_123200_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6385 VSS a_159060_5492# a_159020_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6386 a_104410_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6387 word1.byte2.tinv7.O word1.byte2.tinv6.EN a_124680_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6388 word2.byte2.tinv7.O buf_out13.inv0.I a_113880_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6389 a_150700_11064# a_151030_11904# a_150930_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6390 a_151820_9598# a_151030_9548# a_151650_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6391 VSS a_15780_6952# word5.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6392 VSS buf_out9.inv0.O buf_out9.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6393 a_46020_7976# word6.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6394 a_17220_306# buf_out28.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6395 VSS a_110280_11112# a_111840_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6396 VDD a_157900_9548# a_156900_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6397 a_3820_3276# a_4150_3276# a_4050_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6398 VSS word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6399 Do27_buf buf_out28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6400 word4.byte4.cgate0.inv1.I word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6401 VSS a_15780_3816# word3.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6402 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6403 word8.byte2.cgate0.inv1.I word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6404 a_36120_10500# word7.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6405 a_160500_7976# word6.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6406 a_166260_8628# a_166050_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6407 a_550_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6408 word4.byte4.dff_2.O word4.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6409 a_65350_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6410 a_92280_306# word1.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6411 word2.byte4.cgate0.inv1.I word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6412 VDD buf_out26.inv0.I buf_out26.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X6413 VSS word8.byte1.cgate0.nand0.B a_33420_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6414 word7.byte2.dff_3.O word7.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6415 VDD a_47020_6412# a_46020_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6416 a_62260_9048# a_60420_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6417 a_550_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6418 VSS a_142500_6578# a_144060_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6419 word1.byte4.inv_and.O word1.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6420 word2.byte3.cgate0.inv1.I word2.byte3.cgate0.nand0.A a_73020_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6421 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6422 VSS word1.byte4.tinv2.I a_10020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6423 a_122640_1090# a_122410_140# a_122080_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6424 VDD a_47020_3276# a_46020_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6425 VSS a_142500_3442# a_144060_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6426 a_139900_4792# word4.byte1.dff_7.CLK a_140130_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6427 VSS a_162660_8628# word6.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6428 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6429 buf_sel6.inv1.O buf_sel6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6430 VDD word8.byte1.tinv0.I a_142500_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6431 word7.byte2.cgate0.inv1.I word7.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6432 a_114880_1656# a_115210_2496# a_115110_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6433 a_62580_8628# a_62370_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6434 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6435 a_18780_5912# word4.byte4.cgate0.inv1.O a_18220_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6436 a_139900_1656# word2.byte1.dff_7.CLK a_140130_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6437 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6438 a_56820_6578# buf_out20.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6439 a_11250_5912# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6440 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6441 VDD a_4980_6952# word5.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6442 a_118480_6412# a_118810_6412# a_118710_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6443 a_20820_306# word1.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6444 word3.byte3.tinv7.O word3.byte3.tinv7.EN a_67620_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6445 a_56820_3442# buf_out20.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6446 VSS word5.byte1.cgate0.nand0.B word5.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6447 VSS a_111280_6412# a_110280_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6448 VDD word4.byte4.tinv6.I a_24420_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6449 VSS a_166260_2356# a_166220_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6450 word1.byte1.nand.B word1.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6451 a_111610_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6452 VDD a_4980_3816# word3.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6453 buf_in32.inv1.O buf_in32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6454 a_113880_11112# word8.byte2.tinv3.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6455 a_118480_3276# a_118810_3276# a_118710_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6456 VDD buf_in10.inv0.O buf_in10.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6457 VDD word6.byte3.nand.OUT word6.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6458 VDD a_13620_306# a_15180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6459 VDD a_165100_140# a_164100_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6460 VSS a_111280_3276# a_110280_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6461 VDD word2.byte4.tinv6.I a_24420_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6462 VSS buf_in1.inv0.O buf_in1.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6463 word7.byte1.tinv7.O buf_out1.inv0.I a_167700_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6464 VDD a_26580_5492# a_26540_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6465 buf_in23.inv0.O Di22 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6466 a_113880_1704# word2.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6467 a_4770_1706# word2.byte4.cgate0.inv1.O a_4660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6468 a_154300_140# word1.byte1.dff_7.CLK a_154530_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6469 buf_in30.inv1.O buf_in30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6470 a_19340_9598# a_18550_9548# a_19170_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6471 VSS a_124680_7976# a_126240_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6472 a_58940_12184# a_58150_11904# a_58770_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6473 VSS word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6474 word1.byte1.dff_0.O word1.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6475 VDD a_26580_2356# a_26540_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6476 a_166050_4842# a_165430_5632# a_165940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6477 buf_sel4.inv0.O buf_sel4.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6478 word8.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6479 a_158740_9598# a_156900_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6480 VSS a_47020_7928# a_46020_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6481 a_165330_7978# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6482 VSS a_58980_10088# a_58940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6483 word7.byte2.tinv7.O word7.byte2.tinv0.EN a_103080_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6484 a_166050_1706# a_165430_2496# a_165940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6485 a_95160_9714# word7.byte2.cgate0.nand0.A word7.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6486 a_15780_10088# a_15570_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6487 a_15180_7362# a_14950_6412# a_14620_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6488 a_71760_12850# dec8.and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6489 word6.byte1.dff_0.O word6.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6490 a_65580_12184# word8.byte3.cgate0.inv1.O a_65020_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6491 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6492 a_51180_5912# word4.byte3.cgate0.inv1.O a_50620_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6493 a_162340_10498# a_160500_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6494 VDD word6.byte2.tinv1.I a_106680_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6495 buf_sel7.inv1.O buf_sel7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6496 VDD word5.byte1.nand.B word5.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6497 a_8540_6462# a_7750_6412# a_8370_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6498 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6499 a_15180_4226# a_14950_3276# a_14620_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6500 buf_out14.inv1.O buf_out14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6501 word5.byte4.tinv7.O buf_out28.inv0.I a_17220_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6502 a_25980_2776# word2.byte4.cgate0.inv1.O a_25420_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6503 VDD a_53220_6578# a_54780_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6504 VDD word1.byte1.cgate0.nand0.B word1.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6505 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6506 a_7750_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6507 a_50620_7928# a_50950_8768# a_50850_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6508 a_780_1090# a_550_140# a_220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6509 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6510 VSS buf_in13.inv0.O buf_in13.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6511 a_47020_11064# a_47350_11904# a_47250_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6512 VDD a_161500_11064# a_160500_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6513 a_55170_190# word1.byte3.cgate0.inv1.O a_55060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6514 VDD word3.byte1.nand.B word3.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6515 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6516 VDD a_108840_8628# a_108800_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6517 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6518 a_8540_3326# a_7750_3276# a_8370_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6519 word3.byte4.tinv7.O buf_out28.inv0.I a_17220_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6520 a_58770_11114# a_58150_11904# a_58660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6521 a_151260_9598# word7.byte1.dff_7.CLK a_150700_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6522 VDD a_107680_7928# a_106680_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6523 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6524 VDD a_53220_3442# a_54780_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6525 VDD buf_in16.inv0.O buf_in16.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6526 a_51570_9598# word7.byte3.cgate0.inv1.O a_51460_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6527 a_22050_6462# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6528 a_123200_12184# a_122410_11904# a_123030_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6529 word7.byte3.dff_6.O word7.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6530 VSS buf_in7.inv0.O buf_in7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6531 a_1060_6462# a_120_6462# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6532 VDD buf_in24.inv0.O buf_in24.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6533 VSS word8.byte4.tinv6.I a_24420_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6534 a_22050_3326# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6535 word4.byte4.tinv7.O word4.byte4.tinv0.EN a_2820_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6536 VSS a_165100_1656# a_164100_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6537 word1.byte1.dff_7.O word1.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6538 a_147430_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6539 a_146100_1704# word2.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6540 VSS a_51780_11764# a_51740_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6541 VDD word7.byte3.nand.OUT word7.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6542 a_118480_9548# word7.byte2.dff_7.CLK a_118710_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6543 VSS Di21 buf_in22.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6544 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6545 a_6420_6578# word5.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6546 a_1060_3326# a_120_3326# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6547 VSS word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6548 buf_in22.inv1.O buf_in22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6549 a_147430_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6550 a_144620_4842# word4.byte1.dff_7.CLK a_144450_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6551 word8.byte3.tinv7.O word8.byte3.tinv2.EN a_49620_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6552 word1.byte3.dff_1.O word1.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6553 word6.byte2.dff_3.O word6.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6554 VDD a_166260_8628# word6.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6555 VSS word2.byte4.cgate0.nand0.A a_35760_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6556 VSS word4.byte1.cgate0.nand0.B word4.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6557 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6558 VDD word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6559 a_119600_2776# a_118810_2496# a_119430_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6560 VSS buf_sel2.inv0.I buf_sel2.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6561 a_105240_11764# a_105030_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6562 a_132960_11112# word8.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6563 VSS a_8580_10088# word7.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6564 a_6420_3442# word3.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6565 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6566 a_144620_1706# word2.byte1.dff_7.CLK a_144450_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6567 a_128280_3442# word3.byte2.tinv7.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6568 VSS a_54220_4792# a_53220_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6569 word5.byte2.tinv7.O word5.byte2.tinv2.EN a_110280_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6570 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6571 VDD a_111280_9548# a_110280_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6572 VSS word7.byte4.tinv3.I a_13620_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6573 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6574 VDD word4.buf_sel0.O word4.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6575 word8.byte3.tinv7.O buf_out18.inv0.I a_64020_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6576 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6577 word5.byte3.tinv7.O buf_out22.inv0.I a_49620_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6578 VDD word2.buf_sel0.O word2.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6579 VDD buf_out13.inv0.O buf_out13.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6580 word3.byte3.tinv7.O buf_out22.inv0.I a_49620_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6581 a_28020_7976# buf_out25.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6582 a_18550_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6583 a_61980_6462# word5.byte3.cgate0.inv1.O a_61420_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6584 a_122080_140# a_122410_140# a_122310_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6585 VSS buf_out4.inv0.O Do3_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6586 VSS buf_out25.inv0.I buf_out25.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X6587 VSS a_11020_9548# a_10020_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6588 VDD a_3820_9548# a_2820_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6589 a_142500_7976# word6.byte1.tinv0.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6590 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6591 a_159020_1090# word1.byte1.dff_7.CLK a_158850_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6592 a_61980_3326# word3.byte3.cgate0.inv1.O a_61420_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6593 VDD a_24420_4840# a_25980_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6594 VDD buf_in29.inv0.O buf_in29.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6595 a_26540_11114# word8.byte4.cgate0.inv1.O a_26370_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6596 a_92280_8932# word6.byte2.cgate0.latch0.I0.O word6.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6597 VDD word8.byte2.tinv0.I a_103080_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6598 word1.byte3.tinv7.O word1.byte3.tinv4.EN a_56820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6599 VSS word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6600 VDD a_24420_1704# a_25980_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6601 a_165100_4792# word4.byte1.dff_7.CLK a_165330_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6602 VSS word8.byte3.buf_RE0.O word8.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6603 VSS word3.byte1.inv_and.O a_131700_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6604 VSS a_43420_11064# a_42420_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6605 a_116040_6952# a_115830_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6606 a_165100_1656# word2.byte1.dff_7.CLK a_165330_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6607 VSS a_56820_9714# a_58380_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6608 word4.byte4.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6609 a_25750_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6610 VSS word5.byte1.cgate0.nand0.B word5.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6611 a_126010_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6612 a_123200_9048# a_122410_8768# a_123030_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6613 a_116040_3816# a_115830_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6614 word3.byte2.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B a_93540_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6615 a_54220_7928# word6.byte3.cgate0.inv1.O a_54450_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6616 a_46020_306# word1.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6617 a_161830_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6618 VSS a_144660_5492# a_144620_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6619 word5.byte1.tinv7.O word5.byte1.tinv0.EN a_142500_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6620 word6.byte2.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6621 word7.byte2.tinv7.O buf_out16.inv0.I a_103080_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6622 VSS buf_in16.inv0.O buf_in16.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6623 a_39180_3442# buf_we1.inv1.O word3.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6624 VDD word4.byte3.tinv2.I a_49620_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6625 VSS word5.byte4.tinv5.I a_20820_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6626 a_126010_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6627 VDD a_57820_11064# a_56820_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6628 VDD buf_in9.inv0.O buf_in9.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6629 a_161830_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6630 a_151860_680# a_151650_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6631 a_60420_7976# buf_out19.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6632 VDD word2.byte3.tinv2.I a_49620_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6633 word6.byte1.cgate0.nand0.A word6.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6634 VSS a_139800_190# a_140460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6635 a_50950_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6636 VDD buf_in3.inv0.O buf_in3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6637 VSS a_13620_11112# a_15180_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6638 buf_in26.inv0.O Di25 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6639 word6.byte2.cgate0.inv1.I word6.byte2.cgate0.nand0.A a_95160_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6640 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6641 a_149700_4840# word4.byte1.tinv2.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6642 dec8.and4_1.nand1.OUT dec8.and4_3.nand1.A a_66360_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6643 Do2_buf buf_out3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6644 a_67620_10500# buf_out17.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6645 VSS word6.byte3.tinv3.I a_53220_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6646 a_10020_3442# word3.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6647 VDD Di17 buf_in18.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6648 VDD word5.byte1.tinv3.I a_153300_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6649 word7.byte2.tinv7.O word7.byte2.tinv7.EN a_128280_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6650 a_144060_4842# a_143830_5632# a_143500_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6651 a_100480_1656# a_100810_2496# a_100710_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6652 buf_we3.inv1.O buf_we3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6653 a_7750_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6654 a_110280_6578# buf_out14.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6655 a_44370_4842# a_43750_5632# a_44260_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6656 a_78780_9714# buf_we2.inv1.O word7.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6657 word6.byte1.dff_7.O word6.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6658 VSS word7.byte2.nand.OUT word7.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6659 a_164100_3442# word3.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6660 VDD word3.byte1.tinv3.I a_153300_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6661 word4.byte3.dff_4.O word4.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6662 buf_sel1.inv1.O buf_sel1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6663 a_58770_9598# a_58150_9548# a_58660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6664 VDD a_141060_6952# a_141020_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6665 a_144060_1706# a_143830_2496# a_143500_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6666 a_36120_9714# word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6667 a_44370_1706# a_43750_2496# a_44260_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6668 a_110280_3442# buf_out14.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6669 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.latch0.I0.ENB a_131700_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6670 word5.gt_re3.I word5.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6671 a_43650_2776# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6672 a_112120_190# a_110280_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6673 a_143500_11064# a_143830_11904# a_143730_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6674 word2.byte3.dff_4.O word2.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6675 word3.byte3.tinv7.O word3.byte3.tinv3.EN a_53220_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6676 VSS buf_in15.inv0.O buf_in15.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6677 VDD word1.byte3.nand.OUT word1.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6678 VDD a_141060_3816# a_141020_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6679 word4.gt_re0.OUT buf_sel4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6680 VSS a_151860_2356# a_151820_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6681 a_14850_9048# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6682 a_115110_6462# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6683 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.latch0.I0.ENB a_131700_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6684 a_53220_6578# word5.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6685 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6686 VSS a_164100_306# a_165660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6687 VDD a_150700_140# a_149700_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6688 a_13620_9714# word7.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6689 word2.gt_re0.OUT buf_sel2.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6690 VSS buf_in29.inv0.O buf_in29.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6691 a_112120_5912# a_110280_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6692 word6.byte4.tinv7.O buf_out27.inv0.I a_20820_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6693 a_104640_6462# word5.byte2.dff_7.CLK a_104080_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6694 a_19060_1090# a_17220_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6695 a_115110_3326# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6696 a_220_1656# a_550_2496# a_450_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6697 a_780_12184# word8.byte4.cgate0.inv1.O a_220_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6698 VSS word8.byte1.tinv1.I a_146100_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6699 a_115830_6462# a_115210_6412# a_115720_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6700 VSS a_110280_7976# a_111840_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6701 VDD a_119640_680# word1.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6702 a_104640_3326# word3.byte2.dff_7.CLK a_104080_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6703 a_158460_1090# a_158230_140# a_157900_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6704 buf_in21.inv1.O buf_in21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6705 a_58770_190# a_58150_140# a_58660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6706 a_3820_4792# a_4150_5632# a_4050_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6707 a_118710_190# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6708 a_115830_3326# a_115210_3276# a_115720_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6709 VSS a_112440_10088# a_112400_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6710 a_68700_13636# dec8.and4_2.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6711 buf_in2.inv1.O buf_in2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6712 a_162660_680# a_162450_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6713 VSS a_15780_5492# word4.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6714 a_150930_7978# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6715 a_13620_7976# word6.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6716 a_19380_8628# a_19170_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6717 a_160500_9714# word7.byte1.tinv5.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6718 a_7750_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6719 VDD word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6720 VDD word1.byte2.tinv1.I a_106680_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6721 VSS word4.byte3.tinv5.I a_60420_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6722 a_24420_11112# buf_out26.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6723 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6724 a_108840_680# a_108630_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6725 a_550_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6726 a_17220_4840# word4.byte4.tinv4.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6727 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6728 VSS a_147100_6412# a_146100_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6729 a_58940_7978# word6.byte3.cgate0.inv1.O a_58770_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6730 VDD word5.byte3.cgate0.nand0.A a_75360_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6731 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6732 VDD word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6733 VSS word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6734 VSS buf_out12.inv0.O buf_out12.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6735 a_58660_7362# a_56820_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6736 VSS a_142500_4840# a_144060_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6737 a_54780_9048# word6.byte3.cgate0.inv1.O a_54220_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6738 VSS a_147100_3276# a_146100_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6739 VDD word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6740 VDD word3.byte3.cgate0.nand0.A a_75360_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6741 VDD a_61420_4792# a_60420_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6742 a_42420_4840# word4.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6743 a_26540_10498# word7.byte4.cgate0.inv1.O a_26370_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6744 VSS word1.byte2.tinv2.I a_110280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6745 a_58660_4226# a_56820_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6746 VDD a_159060_6952# word5.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6747 a_167700_8932# word6.byte1.tinv7.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6748 VDD a_61420_1656# a_60420_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6749 a_58980_6952# a_58770_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6750 a_42420_1704# word2.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6751 a_6420_1704# word2.byte4.tinv1.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6752 a_162660_5492# a_162450_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6753 VDD buf_out29.inv0.O Do28_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6754 a_148220_11114# word8.byte1.dff_7.CLK a_148050_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6755 a_25420_9548# a_25750_9548# a_25650_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6756 a_51460_7978# a_49620_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6757 VSS a_150700_1656# a_149700_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6758 a_131700_2660# word2.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6759 VDD a_159060_3816# word3.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6760 VSS buf_out32.inv0.O Do31_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6761 buf_in5.inv1.O buf_in5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6762 Do17_buf buf_out18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6763 VSS a_19380_2356# a_19340_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6764 a_162660_2356# a_162450_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6765 a_58980_3816# a_58770_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6766 a_75720_8932# word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6767 VDD a_12180_6952# word5.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6768 a_118480_4792# a_118810_5632# a_118710_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6769 VSS word2.buf_ck1.I word2.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6770 VSS word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6771 a_108840_8628# a_108630_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6772 a_122920_6462# a_121080_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6773 VDD a_151860_8628# word6.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6774 VDD a_18220_140# a_17220_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6775 a_93540_2660# word2.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6776 VSS a_165100_11064# a_164100_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6777 a_51780_8628# a_51570_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X6778 a_158850_1706# word2.byte1.dff_7.CLK a_158740_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6779 VDD a_12180_3816# word3.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X6780 buf_sel4.inv1.O buf_sel4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6781 VSS a_22980_2356# word2.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6782 a_54220_140# a_54550_140# a_54450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6783 a_113880_3442# word3.byte2.tinv3.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6784 a_147430_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6785 a_122920_3326# a_121080_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6786 a_20820_4840# word4.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6787 VSS word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6788 a_115720_11114# a_113880_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6789 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6790 buf_sel5.inv0.I dec8.and4_4.nand1.OUT a_72300_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6791 VSS a_66180_8628# word6.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6792 word5.byte1.tinv7.O word5.byte1.tinv7.EN a_167700_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6793 a_124680_7976# word6.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6794 VSS word5.byte2.tinv3.I a_113880_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6795 a_155420_190# a_154630_140# a_155250_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6796 a_75720_3442# word3.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6797 a_28020_1092# buf_out25.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6798 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6799 a_18450_7978# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6800 VDD word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6801 word6.byte3.cgate0.nand0.A word6.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6802 a_50850_12184# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6803 VSS word3.byte1.cgate0.nand0.B a_33420_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6804 VDD buf_in11.inv0.O buf_in11.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6805 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6806 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6807 VSS a_149700_1704# a_151260_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6808 a_116000_12184# a_115210_11904# a_115830_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6809 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6810 a_15570_6462# word5.byte4.cgate0.inv1.O a_15460_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6811 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6812 a_119430_9598# word7.byte2.dff_7.CLK a_119320_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6813 word1.byte4.tinv7.O word1.byte4.tinv1.EN a_6420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6814 buf_out11.inv1.O buf_out11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6815 buf_in25.inv0.O Di24 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6816 word5.byte4.dff_7.O word5.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6817 VDD buf_in25.inv0.O buf_in25.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6818 buf_in7.inv0.O Di6 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6819 VSS a_39820_11064# a_39720_11114# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6820 a_50620_11064# word8.byte3.cgate0.inv1.O a_50850_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6821 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6822 VDD a_113880_7976# a_115440_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6823 VDD a_10020_4840# a_11580_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6824 VDD a_57820_6412# a_56820_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6825 a_15570_3326# word3.byte4.cgate0.inv1.O a_15460_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6826 VSS a_153300_6578# a_154860_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6827 VDD a_141060_11764# a_141020_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6828 a_164100_9714# buf_out2.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6829 VSS Di23 buf_in24.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6830 a_114880_6412# word5.byte2.dff_7.CLK a_115110_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6831 word3.byte4.dff_7.O word3.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6832 a_8540_5912# a_7750_5632# a_8370_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6833 a_7650_4842# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6834 VSS word2.gt_re1.O word2.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6835 word6.byte2.inv_and.O word6.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6836 VDD a_10020_1704# a_11580_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6837 VDD a_57820_3276# a_56820_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6838 VDD buf_in31.inv0.O buf_in31.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6839 buf_in17.inv1.O buf_in17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6840 VSS a_153300_3442# a_154860_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6841 word8.byte3.tinv7.O word8.byte3.tinv7.EN a_67620_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6842 word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.latch0.I0.O a_36120_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6843 VSS word2.byte4.buf_RE0.O word2.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6844 a_114880_3276# word3.byte2.dff_7.CLK a_115110_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6845 VDD word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6846 a_7650_1706# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X6847 VSS buf_out17.inv0.O Do16_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6848 a_155140_6462# a_153300_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6849 a_104080_11064# a_104410_11904# a_104310_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6850 VDD word6.byte4.dff_0.O_bar a_2820_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6851 VSS a_55380_6952# a_55340_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6852 VSS word4.byte1.cgate0.nand0.B a_95160_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6853 a_22050_5912# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6854 buf_sel2.inv1.O buf_sel2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6855 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6856 a_39820_140# word1.byte3.cgate0.inv1.O a_40050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6857 a_111610_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6858 word1.byte2.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6859 VSS a_18220_1656# a_17220_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6860 VDD a_166260_6952# a_166220_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6861 VSS word7.byte1.cgate0.nand0.B a_73020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6862 a_162450_7978# word6.byte1.dff_7.CLK a_162340_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6863 VSS word1.byte1.cgate0.nand0.B a_33420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6864 VDD word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6865 word8.byte1.dff_4.O word8.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6866 a_155140_3326# a_153300_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6867 word4.byte1.tinv7.O buf_out4.inv0.I a_156900_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6868 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6869 VDD word4.byte2.tinv0.I a_103080_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6870 VSS a_55380_3816# a_55340_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6871 a_1060_5912# a_120_4842# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6872 VSS word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6873 VDD a_4980_8628# a_4940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6874 VSS a_17220_306# a_18780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6875 a_126240_2776# word2.byte2.dff_7.CLK a_125680_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6876 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6877 a_58380_7978# a_58150_8768# a_57820_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6878 VDD a_166260_3816# a_166220_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6879 a_111610_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6880 a_147430_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6881 a_40050_9048# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6882 a_60420_306# buf_out19.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6883 word7.byte2.dff_2.O word7.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6884 word2.byte1.tinv7.O buf_out4.inv0.I a_156900_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6885 a_4770_6462# a_4150_6412# a_4660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6886 a_25650_190# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6887 VDD word2.byte2.tinv0.I a_103080_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6888 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6889 word6.byte1.nand.B word6.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6890 VDD a_105240_5492# a_105200_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6891 a_131700_306# word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6892 VDD word7.byte1.cgate0.nand0.A word7.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6893 VDD a_104080_4792# a_103080_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6894 word6.byte3.tinv7.O buf_out23.inv0.I a_46020_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6895 a_4770_3326# a_4150_3276# a_4660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6896 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6897 VDD a_105240_2356# a_105200_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6898 VDD buf_out4.inv0.I buf_out4.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X6899 a_15780_680# a_15570_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6900 VDD a_104080_1656# a_103080_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X6901 word6.byte1.tinv7.O word6.byte1.tinv5.EN a_160500_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6902 a_58660_190# a_56820_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6903 buf_in1.inv1.O buf_in1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6904 VSS word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6905 VSS a_57820_7928# a_56820_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6906 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6907 word8.byte2.tinv7.O buf_out11.inv0.I a_121080_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6908 a_25980_7362# a_25750_6412# a_25420_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6909 VDD word5.byte1.buf_RE1.I word5.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6910 a_25980_11114# a_25750_11904# a_25420_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6911 word6.byte1.dff_3.O word6.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6912 VSS word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6913 a_61980_5912# word4.byte3.cgate0.inv1.O a_61420_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6914 a_157900_1656# a_158230_2496# a_158130_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6915 word4.byte3.dff_0.O word4.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6916 VDD A1 dec8.and4_5.nand1.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6917 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6918 VDD word3.byte1.buf_RE1.I word3.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6919 a_25980_4226# a_25750_3276# a_25420_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6920 a_22660_9598# a_20820_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6921 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6922 VDD word8.byte4.tinv1.I a_6420_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6923 VDD a_119640_680# a_119600_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6924 VSS buf_in11.inv0.O buf_in11.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6925 word2.byte3.dff_0.O word2.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6926 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6927 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6928 VSS a_105240_680# a_105200_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6929 a_18220_4792# word4.byte4.cgate0.inv1.O a_18450_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6930 a_100710_6462# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6931 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6932 a_67620_4840# word4.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6933 a_22980_10088# a_22770_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6934 a_148220_10498# word7.byte1.dff_7.CLK a_148050_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6935 word1.byte4.tinv7.O buf_out27.inv0.I a_20820_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6936 a_156900_306# word1.byte1.tinv4.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X6937 a_154630_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6938 a_54550_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6939 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6940 a_18220_1656# word2.byte4.cgate0.inv1.O a_18450_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6941 VSS word5.byte4.nand.OUT word5.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6942 buf_in13.inv1.O buf_in13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6943 a_24420_4840# buf_out26.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6944 VSS buf_out28.inv0.O Do27_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6945 a_100710_3326# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6946 a_67620_1704# word2.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6947 a_116040_5492# a_115830_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X6948 a_14950_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6949 a_156900_1704# word2.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6950 a_24420_1704# buf_out26.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6951 a_62540_9598# a_61750_9548# a_62370_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6952 a_119600_7362# word5.byte2.dff_7.CLK a_119430_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6953 a_115720_9048# a_113880_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X6954 word1.byte2.dff_6.O word1.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6955 a_62260_11114# a_60420_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6956 word2.byte2.tinv7.O word2.byte2.tinv3.EN a_113880_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6957 a_14950_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X6958 a_108010_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6959 a_115720_10498# a_113880_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6960 buf_in24.inv1.O buf_in24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6961 VSS word7.byte1.cgate0.nand0.B a_134580_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6962 VSS word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6963 a_119600_4226# word3.byte2.dff_7.CLK a_119430_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6964 VDD word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6965 a_115210_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6966 a_450_6462# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6967 word7.byte3.inv_and.O word7.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X6968 buf_sel7.inv0.I dec8.and4_6.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6969 VDD a_42420_11112# a_43980_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6970 word7.byte1.tinv7.O word7.byte1.tinv1.EN a_146100_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6971 a_7420_7928# a_7750_8768# a_7650_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X6972 VSS word1.byte3.dff_0.O_bar a_42420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X6973 a_46020_4840# word4.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6974 dec8.and4_6.nand0.OUT dec8.and4_6.nand0.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6975 a_44540_1090# word1.byte3.cgate0.inv1.O a_44370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6976 a_112400_7978# word6.byte2.dff_7.CLK a_112230_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X6977 VSS word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6978 a_33420_2660# word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6979 a_450_3326# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X6980 VSS word5.byte1.buf_RE1.I word5.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6981 a_8370_9598# word7.byte4.cgate0.inv1.O a_8260_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6982 VDD word6.byte1.tinv2.I a_149700_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6983 VDD word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6984 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6985 a_106680_7976# buf_out15.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6986 a_166050_11114# a_165430_11904# a_165940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6987 word2.byte3.dff_2.O word2.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X6988 VDD a_2820_7976# a_4380_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6989 VSS a_101640_6952# word5.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X6990 a_44370_11114# word8.byte3.cgate0.inv1.O a_44260_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6991 a_50620_9548# word7.byte3.cgate0.inv1.O a_50850_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X6992 a_124680_9714# buf_out10.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X6993 VDD a_141060_10088# a_141020_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X6994 a_17220_3442# word3.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X6995 VSS buf_we1.inv0.O buf_we1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X6996 VSS a_21820_9548# a_20820_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X6997 VDD word6.byte3.buf_RE0.O word6.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X6998 a_62370_190# word1.byte3.cgate0.inv1.O a_62260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X6999 VSS a_146100_7976# a_147660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7000 VSS a_101640_3816# word3.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7001 word8.byte3.dff_6.O word8.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7002 VDD buf_in6.inv0.O buf_in6.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7003 a_1060_12184# a_120_11114# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7004 VDD buf_in27.inv0.O buf_in27.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7005 a_62580_11764# a_62370_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7006 word8.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7007 a_123240_2356# a_123030_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7008 a_3820_140# a_4150_140# a_4050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7009 VSS buf_in30.inv0.O buf_in30.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7010 VDD a_50620_9548# a_49620_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7011 word8.byte1.tinv7.O word8.byte1.tinv6.EN a_164100_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7012 a_73020_8932# word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7013 VSS a_48180_8628# a_48140_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7014 word8.byte2.dff_4.O word8.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7015 a_115110_5912# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7016 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7017 VSS buf_sel4.inv0.I buf_sel4.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7018 word6.byte1.dff_4.O word6.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7019 word5.byte4.tinv7.O buf_out31.inv0.I a_6420_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7020 VSS word1.byte3.tinv7.I a_67620_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7021 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7022 VSS word2.byte4.tinv6.I a_24420_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7023 a_65020_140# word1.byte3.cgate0.inv1.O a_65250_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7024 a_124680_306# word1.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7025 a_104640_5912# word4.byte2.dff_7.CLK a_104080_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7026 VSS a_51780_8628# word6.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7027 VSS word4.byte3.nand.OUT word4.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7028 word5.byte1.tinv7.O word5.byte1.tinv3.EN a_153300_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7029 word7.byte2.inv_and.O word7.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7030 VDD word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7031 word3.byte4.tinv7.O buf_out31.inv0.I a_6420_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7032 VDD word4.byte2.tinv7.I a_128280_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7033 VDD word5.byte3.buf_RE0.O word5.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7034 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7035 word1.byte3.cgate0.nand0.A word1.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7036 a_56820_9714# word7.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7037 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7038 a_19060_11114# a_17220_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7039 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7040 a_13620_9714# word7.byte4.tinv3.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7041 VDD word2.byte2.tinv7.I a_128280_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7042 word8.byte4.dff_0.O word8.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7043 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7044 VDD word3.byte3.buf_RE0.O word3.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7045 VDD word8.byte3.inv_and.O a_75720_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7046 a_61750_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7047 VSS a_159060_680# word1.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7048 VDD word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7049 a_105030_9598# word7.byte2.dff_7.CLK a_104920_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7050 VDD a_100380_190# a_101040_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7051 buf_in9.inv1.O buf_in9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7052 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7053 word8.byte1.cgate0.inv1.I word8.byte1.cgate0.nand0.A a_134580_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7054 a_12140_12184# a_11350_11904# a_11970_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7055 buf_in24.inv1.O buf_in24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7056 a_25980_10498# a_25750_9548# a_25420_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7057 a_119320_7978# a_117480_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7058 a_100480_6412# word5.byte2.dff_7.CLK a_100710_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7059 a_15460_4842# a_13620_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7060 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7061 VSS word4.byte2.tinv1.I a_106680_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7062 buf_in5.inv1.O buf_in5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7063 VSS a_12180_680# a_12140_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7064 VDD word1.byte4.dff_0.O_bar a_2820_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7065 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7066 a_15460_1706# a_13620_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7067 a_100480_3276# word3.byte2.dff_7.CLK a_100710_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7068 VSS a_157900_11064# a_156900_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7069 a_154860_4842# a_154630_5632# a_154300_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7070 a_147660_11114# a_147430_11904# a_147100_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7071 word7.byte3.tinv7.O buf_out19.inv0.I a_60420_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7072 a_121080_6578# buf_out11.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7073 a_66360_12850# dec8.and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7074 a_43650_7362# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7075 a_140740_6462# a_139800_6462# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7076 VSS a_40980_6952# a_40940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7077 word1.byte3.tinv7.O word1.byte3.tinv6.EN a_64020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7078 a_15780_5492# a_15570_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7079 VDD a_1380_11764# word8.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7080 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7081 VDD word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7082 a_159060_6952# a_158850_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7083 VSS word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7084 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7085 a_47860_9598# a_46020_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7086 a_58150_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7087 a_154860_1706# a_154630_2496# a_154300_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7088 a_122310_2776# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7089 VSS a_107680_4792# a_106680_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7090 VDD a_151860_6952# a_151820_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7091 a_131700_3442# word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7092 a_121080_3442# buf_out11.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7093 a_140740_3326# a_139800_3326# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7094 a_43650_4226# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7095 word5.gt_re3.I word5.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7096 VSS buf_sel5.inv0.O buf_sel5.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7097 a_15780_2356# a_15570_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7098 VSS a_40980_3816# a_40940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7099 a_54550_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7100 a_166220_9048# a_165430_8768# a_166050_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7101 a_92280_306# word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7102 a_159060_3816# a_158850_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7103 VDD word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7104 word1.byte1.nand.B word1.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7105 a_111840_2776# word2.byte2.dff_7.CLK a_111280_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7106 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7107 VDD buf_sel5.inv0.O buf_sel5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7108 a_43980_7978# a_43750_8768# a_43420_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7109 VDD a_161500_7928# a_160500_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7110 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7111 VDD a_151860_3816# a_151820_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7112 a_58150_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7113 word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.latch0.I0.ENB a_92280_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7114 a_55340_4842# word4.byte3.cgate0.inv1.O a_55170_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7115 a_142500_7976# word6.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7116 a_140740_12184# a_139800_11114# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7117 a_140130_11114# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7118 a_7750_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7119 a_220_6412# word5.byte4.cgate0.inv1.O a_450_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7120 a_125910_6462# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7121 word3.byte2.cgate0.nand0.A word3.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7122 word3.gt_re3.I word3.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7123 a_64020_6578# word5.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7124 a_8260_190# a_6420_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7125 word1.byte3.tinv7.O buf_out23.inv0.I a_46020_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7126 word4.byte4.inv_and.O word4.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7127 a_48180_10088# a_47970_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7128 word8.byte1.nand.B word8.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7129 a_92280_7976# word6.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7130 VDD word6.byte2.buf_RE1.I word6.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7131 word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.latch0.I0.ENB a_92280_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7132 a_55340_1706# word2.byte3.cgate0.inv1.O a_55170_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7133 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7134 a_122920_5912# a_121080_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7135 buf_in27.inv0.O Di26 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7136 buf_out13.inv1.O buf_out13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7137 a_4660_9048# a_2820_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7138 a_20820_6578# word5.byte4.tinv5.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7139 VSS word1.byte1.nand.B a_39180_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7140 a_125910_3326# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7141 a_220_3276# word3.byte4.cgate0.inv1.O a_450_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7142 a_108010_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7143 a_62260_10498# a_60420_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7144 word2.byte4.inv_and.O word2.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7145 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7146 a_134580_8932# word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7147 VDD a_159060_11764# a_159020_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7148 a_108010_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7149 buf_in29.inv1.O buf_in29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7150 a_4980_8628# a_4770_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7151 a_21820_6412# a_22150_6412# a_22050_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7152 a_161730_1090# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7153 VDD a_42420_9714# a_43980_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7154 VSS word6.gt_re1.O word6.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7155 Do1_buf buf_out2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7156 Do23_buf buf_out24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7157 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7158 VSS word2.buf_sel0.O word2.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7159 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7160 VDD a_139800_11114# a_140460_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7161 a_21820_3276# a_22150_3276# a_22050_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7162 VSS word7.byte2.tinv4.I a_117480_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7163 a_53220_7976# word6.byte3.tinv3.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7164 a_100710_190# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7165 a_166050_9598# a_165430_9548# a_165940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7166 a_143500_1656# a_143830_2496# a_143730_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7167 a_15570_4842# word4.byte4.cgate0.inv1.O a_15460_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7168 a_153300_6578# buf_out5.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7169 VDD buf_out17.inv0.I buf_out17.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X7170 a_126630_11114# a_126010_11904# a_126520_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7171 VSS a_123240_2356# word2.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7172 word7.byte1.nand.OUT buf_we4.inv1.O a_129540_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7173 VDD a_55380_8628# word6.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7174 a_28020_5796# word4.byte4.tinv7.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7175 VSS a_157900_6412# a_156900_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7176 word4.byte4.dff_7.O word4.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7177 a_153300_11112# word8.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7178 a_132960_7976# word6.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7179 word7.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7180 VSS word7.byte1.cgate0.nand0.B word7.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7181 a_90120_306# word1.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7182 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7183 a_153300_3442# buf_out5.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7184 VSS a_153300_4840# a_154860_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7185 VSS a_157900_3276# a_156900_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7186 a_121080_4840# word4.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7187 VDD buf_sel6.inv0.O buf_sel6.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7188 VSS word7.byte4.inv_and.O a_36120_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7189 word7.byte3.dff_6.O word7.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7190 VSS a_126840_6952# word5.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7191 VDD buf_in14.inv0.O buf_in14.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7192 VSS word3.byte3.dff_0.O_bar a_42420_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7193 word5.gt_re3.I word5.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7194 word4.byte1.cgate0.latch0.I0.O word4.byte1.cgate0.latch0.I0.O a_132960_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7195 a_158130_6462# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7196 a_7420_11064# a_7750_11904# a_7650_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7197 VSS a_126840_11764# a_126800_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7198 word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.latch0.I0.O a_36120_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7199 a_121080_1704# word2.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7200 a_10020_4840# buf_out30.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7201 VDD a_19380_6952# a_19340_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7202 a_62260_1090# a_60420_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7203 VSS a_126840_3816# word3.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7204 a_104080_9548# a_104410_9548# a_104310_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7205 a_450_190# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7206 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.latch0.I0.O a_132960_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7207 word8.byte2.tinv7.O word8.byte2.tinv6.EN a_124680_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7208 a_155140_5912# a_153300_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7209 a_158130_3326# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7210 VSS a_55380_5492# a_55340_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7211 VDD word6.byte4.tinv2.I a_10020_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7212 a_10020_1704# buf_out30.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7213 word1.byte4.dff_7.O word1.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7214 VDD a_19380_3816# a_19340_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7215 VSS Di25 buf_in26.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7216 a_158850_6462# a_158230_6412# a_158740_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7217 VDD a_141060_11764# word8.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7218 VDD a_166260_11764# word8.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7219 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7220 VDD a_22980_6952# word5.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7221 VDD a_162660_680# word1.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7222 a_134580_306# word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7223 a_47250_9598# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7224 VDD Di7 buf_in8.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7225 a_62580_680# a_62370_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7226 buf_in20.inv1.O buf_in20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7227 VSS a_19380_11764# word8.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7228 VDD a_12180_8628# a_12140_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7229 a_158850_3326# a_158230_3276# a_158740_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7230 a_100810_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7231 VSS a_155460_10088# a_155420_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7232 Do31_buf buf_out32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7233 VDD a_22980_3816# word3.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7234 word4.byte2.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7235 VSS a_103080_306# a_104640_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7236 VSS word2.byte3.tinv2.I a_49620_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7237 a_125910_190# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7238 a_64020_11112# word8.byte3.tinv6.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7239 VDD word1.byte1.tinv2.I a_149700_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7240 a_19060_10498# a_17220_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7241 word6.byte4.tinv7.O word6.byte4.tinv3.EN a_13620_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7242 a_151650_7978# a_151030_8768# a_151540_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7243 VSS a_39720_6462# a_40380_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7244 VSS word5.byte2.tinv6.I a_124680_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7245 a_60420_4840# word4.byte3.tinv5.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7246 VDD word7.gt_re1.O word7.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7247 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7248 a_106680_306# buf_out15.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7249 VSS buf_sel1.inv0.O buf_sel1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7250 a_22770_1706# word2.byte4.cgate0.inv1.O a_22660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7251 VDD a_149700_6578# a_151260_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7252 word7.byte4.dff_1.O word7.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7253 VDD a_11020_11064# a_10020_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7254 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7255 VDD word5.byte3.tinv6.I a_64020_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7256 a_116040_680# a_115830_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7257 VSS a_39720_3326# a_40380_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7258 VDD a_1380_5492# a_1340_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7259 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7260 VDD word1.byte3.buf_RE0.O word1.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7261 VDD a_149700_3442# a_151260_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7262 VDD word4.byte3.cgate0.nand0.A word4.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7263 a_8260_7978# a_6420_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7264 word5.byte2.dff_1.O word5.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7265 VDD word3.byte3.tinv6.I a_64020_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7266 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7267 buf_we4.inv0.O WE3 VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X7268 word7.byte1.dff_5.O word7.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7269 VDD a_124680_306# a_126240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7270 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7271 VDD a_1380_2356# a_1340_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7272 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7273 VDD word2.byte3.cgate0.nand0.A word2.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7274 buf_in13.inv1.O buf_in13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7275 word4.byte3.tinv7.O buf_out24.inv0.I a_42420_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7276 word3.byte2.dff_1.O word3.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7277 VDD word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7278 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7279 VSS a_111280_11064# a_110280_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7280 VDD word7.byte1.cgate0.nand0.B word7.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7281 VDD word7.byte1.inv_and.O a_131700_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7282 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7283 VDD word7.byte1.tinv4.I a_156900_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7284 buf_in4.inv1.O buf_in4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7285 a_147660_10498# a_147430_9548# a_147100_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7286 a_8580_8628# a_8370_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7287 a_162340_2776# a_160500_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7288 a_26540_6462# a_25750_6412# a_26370_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7289 VSS a_62580_2356# a_62540_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7290 word2.byte3.tinv7.O buf_out24.inv0.I a_42420_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7291 VDD a_1380_10088# word7.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7292 buf_in25.inv1.O buf_in25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7293 VDD a_61420_140# a_60420_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7294 word1.byte1.dff_0.O word1.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7295 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.latch0.I0.O a_131700_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7296 a_26540_3326# a_25750_3276# a_26370_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7297 a_100710_5912# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7298 buf_sel3.inv0.I dec8.and4_2.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7299 a_165940_6462# a_164100_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7300 VDD a_125680_11064# a_124680_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7301 word2.gt_re0.OUT buf_sel2.inv1.O a_82020_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7302 a_126240_7362# a_126010_6412# a_125680_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7303 VDD buf_in19.inv0.O buf_in19.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7304 VDD word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7305 a_50620_140# word1.byte3.cgate0.inv1.O a_50850_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7306 a_140130_10498# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7307 a_101320_12184# a_100380_11114# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7308 a_156900_3442# word3.byte1.tinv4.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7309 VSS a_3820_11064# a_2820_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7310 a_110280_9714# word7.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7311 a_165940_3326# a_164100_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7312 VDD word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7313 buf_sel7.inv0.O buf_sel7.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7314 a_49620_11112# word8.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7315 a_111610_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7316 a_118710_9048# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7317 a_126240_4226# a_126010_3276# a_125680_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7318 a_61420_140# a_61750_140# a_61650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7319 VDD word3.byte2.cgate0.inv1.I word3.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7320 word4.byte4.tinv7.O word4.byte4.tinv5.EN a_20820_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7321 VSS word5.byte1.tinv4.I a_156900_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7322 a_167700_7976# word6.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7323 a_61650_7978# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7324 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7325 word5.byte4.cgate0.nand0.A word5.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7326 word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.latch0.I0.ENB a_75720_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7327 word6.byte2.tinv7.O buf_out10.inv0.I a_124680_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7328 a_24420_6578# word5.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7329 a_162620_190# a_161830_140# a_162450_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7330 VDD a_159060_10088# a_159020_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7331 VDD a_114880_4792# a_113880_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7332 a_46020_6578# word5.byte3.tinv1.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7333 word3.byte3.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7334 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7335 word4.byte4.cgate0.inv1.I word4.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7336 a_108800_9598# a_108010_9548# a_108630_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7337 word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.latch0.I0.ENB a_75720_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7338 a_450_5912# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7339 a_24420_3442# word3.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7340 buf_out10.inv1.O buf_out10.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7341 VSS a_26580_10088# word7.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7342 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7343 VDD a_114880_1656# a_113880_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7344 a_55380_11764# a_55170_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7345 a_108800_190# a_108010_140# a_108630_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7346 word2.byte4.cgate0.inv1.I word2.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7347 Do0_buf buf_out1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7348 a_104920_7978# a_103080_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7349 Do22_buf buf_out23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7350 VDD a_139800_9598# a_140460_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7351 a_47020_6412# a_47350_6412# a_47250_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7352 a_117480_7976# word6.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7353 a_141060_2356# a_140850_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7354 a_157900_6412# word5.byte1.dff_7.CLK a_158130_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7355 buf_in30.inv0.O Di29 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7356 a_126630_9598# a_126010_9548# a_126520_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7357 a_129540_8932# word6.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7358 a_40150_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7359 word8.byte2.dff_2.O word8.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7360 VSS word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7361 a_40660_190# a_39720_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7362 a_47020_3276# a_47350_3276# a_47250_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7363 VSS a_101640_5492# word4.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7364 a_148050_190# word1.byte1.dff_7.CLK a_147940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7365 word4.byte2.dff_5.O word4.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7366 a_11350_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7367 a_157900_3276# word3.byte1.dff_7.CLK a_158130_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7368 VSS a_165100_140# a_164100_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7369 VDD a_39820_4792# a_39720_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7370 a_43750_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7371 VSS a_61420_1656# a_60420_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7372 a_42420_1704# word2.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7373 word2.byte2.dff_5.O word2.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7374 a_142500_306# word1.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7375 a_154630_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7376 a_151820_9048# a_151030_8768# a_151650_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7377 a_150700_7928# word6.byte1.dff_7.CLK a_150930_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7378 a_2820_7976# buf_out32.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7379 a_103080_306# word1.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7380 VDD a_39820_1656# a_39720_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7381 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7382 a_43750_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7383 VDD word4.byte1.tinv1.I a_146100_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7384 a_40940_4842# word4.byte3.cgate0.inv1.O a_40770_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7385 buf_sel8.inv0.O buf_sel8.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7386 word8.byte2.dff_5.O word8.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7387 a_92280_1092# word1.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7388 VDD word1.byte2.buf_RE1.I word1.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7389 a_101640_10088# a_101430_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7390 VSS word1.byte3.buf_RE0.O word1.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7391 VSS word3.byte3.tinv7.I a_67620_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7392 VSS word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7393 a_154630_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7394 VDD word8.byte3.tinv3.I a_53220_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7395 a_119640_11764# a_119430_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7396 VSS word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7397 VDD word2.byte1.tinv1.I a_146100_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7398 a_40940_1706# word2.byte3.cgate0.inv1.O a_40770_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7399 buf_in13.inv1.O buf_in13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7400 VDD a_148260_5492# a_148220_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7401 VDD a_101640_11764# word8.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7402 VDD a_141060_10088# word7.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7403 VDD a_166260_10088# word7.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7404 VDD buf_in16.inv0.I buf_in16.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7405 VSS a_122080_9548# a_121080_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7406 VDD a_148260_2356# a_148220_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7407 VSS Di6 buf_in7.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7408 buf_in24.inv1.O buf_in24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7409 VSS word6.byte3.buf_RE0.O word6.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7410 VSS a_60420_1704# a_61980_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7411 a_82020_8932# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7412 a_22980_680# a_22770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7413 word7.byte3.tinv7.O buf_out21.inv0.I a_53220_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7414 a_65860_190# a_64020_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7415 a_124680_4840# word4.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7416 buf_in31.inv1.O buf_in31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7417 a_123200_1090# word1.byte2.dff_7.CLK a_123030_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7418 VDD a_104080_140# a_103080_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7419 a_11580_12184# word8.byte4.cgate0.inv1.O a_11020_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7420 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7421 VSS word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7422 word4.byte3.cgate0.nand0.A word4.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7423 buf_in22.inv0.O Di21 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7424 word5.byte3.dff_2.O word5.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7425 a_132960_1092# word1.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7426 buf_sel2.inv0.I dec8.and4_1.nand1.OUT a_66900_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7427 VSS a_64020_6578# a_65580_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7428 VDD a_40980_8628# word6.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7429 a_147660_2776# word2.byte1.dff_7.CLK a_147100_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7430 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7431 word8.byte1.cgate0.nand0.A word8.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7432 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7433 VDD word5.byte1.buf_RE1.I word5.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7434 a_47970_1706# word2.byte3.cgate0.inv1.O a_47860_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7435 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7436 VSS buf_sel2.inv0.O buf_sel2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7437 a_128280_306# word1.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7438 a_140130_2776# buf_in8.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7439 word3.byte1.tinv7.O word3.byte1.tinv2.EN a_149700_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7440 VSS word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7441 word3.byte3.dff_2.O word3.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7442 word2.byte3.dff_5.O word2.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7443 VSS a_64020_3442# a_65580_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7444 a_61420_4792# word4.byte3.cgate0.inv1.O a_61650_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7445 word5.byte1.nand.B word5.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7446 word8.gt_re3.I word8.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7447 a_158130_11114# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7448 a_158740_12184# a_156900_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7449 VDD word3.byte1.buf_RE1.I word3.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7450 word4.byte2.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7451 a_61420_1656# word2.byte3.cgate0.inv1.O a_61650_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7452 a_28020_3442# word3.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7453 a_143730_6462# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7454 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7455 a_123240_6952# a_123030_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7456 VSS a_112440_680# a_112400_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7457 word3.byte1.nand.B word3.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7458 a_40150_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7459 a_48140_2776# a_47350_2496# a_47970_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7460 VDD word1.byte4.tinv2.I a_10020_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7461 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7462 a_101430_6462# word5.byte2.dff_7.CLK a_101320_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7463 a_58050_190# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7464 a_95160_306# word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7465 a_140740_5912# a_139800_4842# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7466 a_22980_11764# a_22770_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7467 VDD word6.byte1.cgate0.nand0.B word6.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7468 word4.byte3.tinv7.O buf_out17.inv0.I a_67620_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7469 a_164100_306# word1.byte1.tinv6.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7470 a_143730_3326# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7471 VSS a_40980_5492# a_40940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7472 a_19340_9048# a_18550_8768# a_19170_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7473 a_123240_3816# a_123030_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7474 a_159060_5492# a_158850_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7475 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7476 a_58150_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7477 VDD a_14620_7928# a_13620_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7478 VSS word4.byte4.dff_0.O_bar a_2820_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7479 buf_we1.inv1.O buf_we1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7480 a_101430_3326# word3.byte2.dff_7.CLK a_101320_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7481 word2.byte3.tinv7.O buf_out17.inv0.I a_67620_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7482 buf_in8.inv1.O buf_in8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7483 word8.byte4.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7484 a_131700_12068# word8.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7485 buf_in29.inv1.O buf_in29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7486 a_158740_9048# a_156900_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7487 a_48180_680# a_47970_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7488 word1.byte1.dff_7.O word1.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7489 VSS a_58980_8628# a_58940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7490 word2.byte1.tinv7.O word2.byte1.tinv4.EN a_156900_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7491 VSS word2.byte2.tinv0.I a_103080_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7492 a_125910_5912# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7493 VSS buf_in18.inv0.O buf_in18.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7494 VDD a_156900_11112# a_158460_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7495 a_111610_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7496 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7497 VSS a_220_9548# a_120_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7498 a_158230_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7499 CLK buf_ck.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7500 word4.byte1.nand.B word4.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7501 a_125910_12184# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7502 word8.byte4.tinv7.O buf_out30.inv0.I a_10020_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7503 a_155420_7978# word6.byte1.dff_7.CLK a_155250_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7504 a_14850_1090# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7505 VDD a_3820_4792# a_2820_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7506 a_44260_6462# a_42420_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7507 VSS a_104080_1656# a_103080_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7508 a_15740_190# a_14950_140# a_15570_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7509 word4.byte3.tinv7.O word4.byte3.tinv1.EN a_46020_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7510 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7511 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7512 a_151260_9048# word6.byte1.dff_7.CLK a_150700_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7513 a_151650_11114# word8.byte1.dff_7.CLK a_151540_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7514 VSS word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7515 a_51570_7978# word6.byte3.cgate0.inv1.O a_51460_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7516 word1.byte2.dff_0.O word1.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7517 VDD a_3820_1656# a_2820_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7518 a_49620_6578# word5.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7519 a_40380_4842# a_40150_5632# a_39820_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7520 a_21820_4792# a_22150_5632# a_22050_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7521 a_44260_3326# a_42420_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7522 a_4150_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7523 buf_out16.inv1.O buf_out16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7524 word6.byte3.dff_6.O word6.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7525 VSS a_144660_6952# word5.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7526 a_60420_3442# word3.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7527 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7528 a_44580_6952# a_44370_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7529 VDD a_110280_306# a_111840_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7530 a_40380_1706# a_40150_2496# a_39820_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7531 a_49620_3442# word3.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7532 buf_in9.inv1.O buf_in9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7533 VSS word5.byte4.buf_RE0.O word5.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7534 a_4150_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7535 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7536 VSS a_144660_3816# word3.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7537 VSS a_141060_680# word1.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7538 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7539 VDD word7.byte1.nand.OUT word7.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7540 a_44580_3816# a_44370_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7541 VDD a_159060_11764# word8.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7542 a_166260_2356# a_166050_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7543 Do25_buf buf_out26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7544 VDD Di2 buf_in3.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7545 VSS a_18220_140# a_17220_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7546 a_122310_7362# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7547 a_65350_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7548 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7549 VDD word7.byte3.buf_RE0.O word7.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7550 VSS a_8580_8628# word6.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7551 VSS a_126840_5492# word4.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7552 a_111840_7362# a_111610_6412# a_111280_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7553 a_122310_4226# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7554 a_158130_5912# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7555 word7.byte2.dff_5.O word7.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7556 VDD buf_out18.inv0.O Do17_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7557 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7558 a_67620_2660# word2.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7559 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7560 a_54780_1090# a_54550_140# a_54220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7561 a_167700_1092# word1.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7562 VSS a_106680_6578# a_108240_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7563 a_24420_1704# word2.byte4.tinv6.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7564 a_111840_4226# a_111610_3276# a_111280_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7565 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7566 VSS word5.byte1.tinv0.I a_142500_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7567 VDD a_101640_10088# word7.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7568 a_126840_10088# a_126630_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7569 word1.byte2.tinv7.O buf_out10.inv0.I a_124680_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7570 VDD buf_sel1.inv0.O buf_sel1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7571 word8.byte3.cgate0.nand0.A word8.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7572 VSS word7.byte2.buf_RE1.I word7.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7573 word1.byte2.dff_7.O word1.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7574 VSS a_106680_3442# a_108240_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7575 a_128280_4840# buf_out9.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7576 word6.byte2.tinv7.O buf_out14.inv0.I a_110280_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7577 VSS word5.byte2.inv_and.O a_92280_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7578 word7.byte3.tinv7.O word7.byte3.tinv4.EN a_56820_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7579 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7580 a_118810_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7581 a_148050_9598# word7.byte1.dff_7.CLK a_147940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7582 a_128280_1704# buf_out9.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7583 buf_in15.inv1.O buf_in15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7584 VSS a_43420_6412# a_42420_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7585 VDD a_154300_6412# a_153300_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7586 VDD word7.byte1.tinv2.I a_149700_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7587 a_108840_680# a_108630_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7588 a_118810_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7589 buf_in6.inv1.O buf_in6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7590 a_13620_9714# buf_out29.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7591 VSS a_39720_4842# a_40380_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7592 VSS a_43420_3276# a_42420_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7593 a_121080_11112# word8.byte2.tinv5.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7594 a_28020_12068# word8.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7595 VDD a_154300_3276# a_153300_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7596 a_143500_6412# word5.byte1.dff_7.CLK a_143730_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7597 VDD a_123240_6952# word5.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7598 VSS word4.byte1.tinv2.I a_149700_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7599 word7.byte4.dff_3.O word7.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7600 buf_in21.inv0.O Di20 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7601 VSS a_56820_7976# a_58380_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7602 a_64020_7976# word6.byte3.tinv6.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7603 VDD a_66180_680# word1.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7604 a_143500_3276# word3.byte1.dff_7.CLK a_143730_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7605 a_106680_4840# word4.byte2.tinv1.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7606 VSS a_139800_9598# a_140460_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7607 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7608 VDD a_123240_3816# word3.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7609 word4.byte2.dff_1.O word4.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7610 a_164100_6578# buf_out2.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7611 dec8.and4_3.nand0.OUT A0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7612 a_119320_12184# a_117480_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7613 a_158130_10498# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7614 a_2820_306# buf_out32.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7615 a_71220_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7616 word7.byte3.cgate0.inv1.I word7.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7617 a_165330_2776# buf_in1.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7618 VSS word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7619 a_164100_3442# buf_out2.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7620 VSS word4.byte3.buf_RE0.O word4.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7621 VSS word3.byte2.tinv5.I a_121080_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7622 VDD word4.byte1.inv_and.O a_131700_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7623 VDD buf_sel7.inv0.O buf_sel7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7624 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7625 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7626 a_55170_7978# a_54550_8768# a_55060_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7627 a_26540_5912# a_25750_5632# a_26370_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7628 a_22980_10088# a_22770_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7629 word5.byte4.dff_0.O word5.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7630 a_25650_4842# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7631 word6.byte3.dff_7.O word6.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7632 VDD word6.byte1.cgate0.nand0.B word6.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7633 VDD word5.byte4.buf_RE0.O word5.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7634 VDD word2.byte1.inv_and.O a_131700_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7635 word3.byte3.cgate0.inv1.O word3.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7636 word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.latch0.I0.O a_93540_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7637 word6.byte1.tinv7.O buf_out8.inv0.I a_142500_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7638 a_126630_6462# word5.byte2.dff_7.CLK a_126520_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7639 a_25650_1706# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7640 word3.byte4.dff_0.O word3.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7641 a_165940_5912# a_164100_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7642 word5.byte3.tinv7.O word5.byte3.tinv6.EN a_64020_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7643 VDD buf_we1.inv1.O word4.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7644 a_144660_11764# a_144450_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7645 VSS a_108840_2356# a_108800_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7646 VDD word3.byte4.buf_RE0.O word3.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7647 VDD word6.byte4.tinv5.I a_20820_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7648 word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.latch0.I0.O a_93540_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7649 a_54220_11064# a_54550_11904# a_54450_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7650 a_126630_3326# word3.byte2.dff_7.CLK a_126520_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7651 VDD a_121080_4840# a_122640_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7652 VDD a_156900_9714# a_158460_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7653 a_65970_11114# a_65350_11904# a_65860_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7654 a_58050_9598# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7655 VDD buf_we1.inv1.O word2.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7656 buf_in28.inv1.O buf_in28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7657 a_115440_9598# word7.byte2.dff_7.CLK a_114880_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7658 VDD a_22980_8628# a_22940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7659 VSS a_154300_7928# a_153300_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7660 a_11580_6462# word5.byte4.cgate0.inv1.O a_11020_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7661 a_134580_8932# word6.byte1.cgate0.nand0.A word6.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7662 VSS word2.byte2.tinv7.I a_128280_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7663 VDD a_121080_1704# a_122640_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7664 VSS buf_out18.inv0.I buf_out18.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X7665 VSS buf_in5.inv0.O buf_in5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7666 a_106680_11112# word8.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7667 a_22770_6462# a_22150_6412# a_22660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7668 a_162450_190# a_161830_140# a_162340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7669 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7670 VSS a_44580_680# a_44540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7671 a_11580_3326# word3.byte4.cgate0.inv1.O a_11020_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7672 VDD buf_in22.inv0.O buf_in22.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7673 VSS word1.byte1.nand.OUT word1.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7674 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7675 a_112230_11114# word8.byte2.dff_7.CLK a_112120_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7676 a_22770_3326# a_22150_3276# a_22660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7677 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.latch0.I0.ENB a_131700_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7678 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7679 a_107910_7978# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7680 a_40050_1090# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7681 a_10020_4840# word4.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7682 VDD a_2820_11112# a_4380_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7683 VSS a_166260_2356# word2.byte1.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7684 word2.byte2.dff_3.O word2.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7685 a_117480_9714# word7.byte2.tinv4.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7686 a_7650_190# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7687 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7688 a_10020_1704# word2.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7689 a_47020_4792# a_47350_5632# a_47250_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7690 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7691 VSS word7.buf_ck1.I word7.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7692 a_65580_4842# a_65350_5632# a_65020_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7693 a_112440_11764# a_112230_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7694 VDD word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7695 a_164100_4840# word4.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7696 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7697 a_4940_9598# a_4150_9548# a_4770_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7698 VDD word1.byte1.cgate0.nand0.B word1.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7699 VSS word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7700 a_162340_7362# a_160500_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7701 word5.byte1.cgate0.inv1.I word5.byte1.cgate0.nand0.A a_134580_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7702 VDD a_159060_10088# word7.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7703 word6.gt_re3.I word6.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7704 VDD a_62580_6952# a_62540_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7705 a_65580_1706# a_65350_2496# a_65020_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7706 a_164100_1704# word2.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7707 a_42420_3442# word3.byte3.tinv0.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7708 VDD word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7709 a_4770_11114# word8.byte4.cgate0.inv1.O a_4660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7710 word4.byte3.tinv7.O buf_out21.inv0.I a_53220_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7711 VDD word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7712 a_105200_6462# a_104410_6412# a_105030_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7713 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7714 a_147100_9548# a_147430_9548# a_147330_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7715 VSS a_120_190# a_780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7716 a_162340_4226# a_160500_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7717 a_43750_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7718 VDD a_62580_3816# a_62540_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7719 a_53220_7976# word6.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7720 word2.byte3.tinv7.O buf_out21.inv0.I a_53220_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7721 VDD buf_out11.inv0.O buf_out11.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7722 VSS a_112440_8628# a_112400_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7723 VSS word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7724 a_105200_3326# a_104410_3276# a_105030_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7725 a_101320_4842# a_100380_4842# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7726 Do6_buf buf_out7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7727 word1.byte1.dff_3.O word1.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7728 VSS word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7729 a_162060_190# word1.byte1.dff_7.CLK a_161500_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7730 VSS buf_out2.inv0.O Do1_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7731 VSS buf_out24.inv0.O Do23_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7732 VDD a_139900_7928# a_139800_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7733 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7734 a_101320_1706# a_100380_1706# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7735 word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.latch0.I0.O a_92280_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7736 a_143830_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7737 VSS a_161500_4792# a_160500_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7738 a_142500_4840# word4.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7739 VDD Di30 buf_in31.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7740 buf_in17.inv0.O Di16 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7741 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7742 word2.byte4.inv_and.O word2.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7743 VDD a_120_4842# a_780_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7744 VSS word4.byte2.buf_RE1.I word4.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7745 a_92280_5796# word4.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7746 VDD word8.byte2.tinv2.I a_110280_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7747 VDD a_108840_8628# word6.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7748 a_141020_7978# word6.byte1.dff_7.CLK a_140850_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7749 VSS a_110280_306# a_111840_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7750 VSS word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7751 VSS word5.byte1.tinv7.I a_167700_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7752 VDD a_120_1706# a_780_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7753 VDD buf_sel2.inv0.O buf_sel2.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7754 word5.byte2.cgate0.inv1.I word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7755 a_103080_6578# word5.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7756 VSS word7.gt_re0.OUT word7.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7757 VSS a_50620_11064# a_49620_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7758 a_124680_6578# word5.byte2.tinv6.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7759 a_40380_11114# a_40150_11904# a_39820_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7760 a_147100_140# a_147430_140# a_147330_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7761 a_33420_3442# word3.byte4.cgate0.nand0.A word3.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7762 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7763 buf_in14.inv1.O buf_in14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7764 a_54220_1656# a_54550_2496# a_54450_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7765 a_103080_3442# word3.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7766 word3.byte2.cgate0.inv1.I word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7767 a_58150_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7768 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7769 a_75360_6578# word5.byte1.cgate0.nand0.B word5.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7770 a_123240_680# a_123030_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7771 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7772 word5.byte1.dff_2.O word5.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7773 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7774 a_141060_6952# a_140850_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7775 a_115720_1090# a_113880_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7776 VDD word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7777 VSS word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7778 a_21820_11064# word8.byte4.cgate0.inv1.O a_22050_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7779 a_25420_7928# a_25750_8768# a_25650_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7780 word7.byte2.tinv7.O buf_out14.inv0.I a_110280_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7781 a_40150_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7782 a_125680_6412# a_126010_6412# a_125910_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7783 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7784 VSS a_15780_11764# a_15740_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7785 word3.byte1.dff_2.O word3.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7786 VSS a_64020_4840# a_65580_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7787 a_141060_3816# a_140850_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7788 a_40660_12184# a_39720_11114# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7789 a_149700_11112# word8.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7790 a_26370_9598# word7.byte4.cgate0.inv1.O a_26260_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7791 buf_in3.inv1.O buf_in3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7792 word8.byte4.tinv7.O word8.byte4.tinv3.EN a_13620_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7793 a_50950_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7794 a_125680_3276# a_126010_3276# a_125910_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X7795 a_40150_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7796 a_7420_140# word1.byte4.cgate0.inv1.O a_7650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7797 word1.byte3.dff_5.O word1.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7798 a_132960_5796# word4.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7799 VSS buf_in20.inv0.O buf_in20.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7800 VDD a_20820_7976# a_22380_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7801 a_35760_8932# word6.byte1.cgate0.nand0.B word6.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7802 VSS a_164100_9714# a_165660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7803 a_122410_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7804 a_121080_1704# word2.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7805 VSS a_20820_11112# a_22380_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7806 a_143730_5912# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7807 word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B a_132960_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7808 dec8.and4_5.nand1.OUT A2 a_73560_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7809 word8.byte4.tinv7.O buf_out25.inv0.I a_28020_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7810 a_161500_7928# word6.byte1.dff_7.CLK a_161730_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7811 a_101430_4842# word4.byte2.dff_7.CLK a_101320_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7812 a_122410_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7813 VDD a_100480_4792# a_100380_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7814 a_10020_1704# word2.byte4.tinv2.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7815 a_153300_9714# word7.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7816 a_112440_10088# a_112230_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7817 word1.byte2.tinv7.O buf_out14.inv0.I a_110280_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7818 VSS a_66180_10088# a_66140_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7819 a_144660_10088# a_144450_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7820 VDD a_100480_1656# a_100380_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7821 a_113880_4840# buf_out13.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7822 VSS word4.byte4.tinv2.I a_10020_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7823 VDD a_146100_306# a_147660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7824 a_119430_7978# word6.byte2.dff_7.CLK a_119320_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7825 a_108240_4842# a_108010_5632# a_107680_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7826 word6.byte1.tinv7.O buf_out1.inv0.I a_167700_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7827 VSS word8.buf_ck1.I word8.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7828 VDD word6.byte2.tinv3.I a_113880_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7829 a_65970_9598# a_65350_9548# a_65860_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7830 a_113880_1704# buf_out13.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X7831 word8.byte3.dff_0.O word8.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7832 a_4380_9598# word7.byte4.cgate0.inv1.O a_3820_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7833 a_75720_4840# word4.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7834 word8.byte3.dff_7.O word8.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7835 word5.byte4.tinv7.O buf_out26.inv0.I a_24420_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7836 a_108240_1706# a_108010_2496# a_107680_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7837 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7838 VDD a_60420_6578# a_61980_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7839 VDD word4.byte1.cgate0.nand0.B word4.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7840 buf_in27.inv1.O buf_in27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7841 VSS buf_in13.inv0.O buf_in13.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7842 VDD a_48180_680# a_48140_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7843 VDD a_116040_8628# a_116000_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7844 VSS word6.byte1.tinv5.I a_160500_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7845 a_75720_1704# word2.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7846 word3.byte4.tinv7.O buf_out26.inv0.I a_24420_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7847 a_147940_7978# a_146100_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7848 VDD a_60420_3442# a_61980_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7849 a_44260_5912# a_42420_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7850 VDD a_11020_4792# a_10020_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7851 a_116000_190# a_115210_140# a_115830_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7852 a_20820_9714# word7.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7853 VDD word2.byte1.cgate0.nand0.B word2.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7854 a_147660_7362# a_147430_6412# a_147100_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7855 a_47970_6462# a_47350_6412# a_47860_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7856 VDD a_114880_140# a_113880_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7857 VDD a_2820_9714# a_4380_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7858 word6.byte2.tinv7.O word6.byte2.tinv4.EN a_117480_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7859 a_140130_7362# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7860 VSS word6.byte1.nand.OUT word6.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7861 VDD a_51780_680# word1.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7862 VDD a_11020_1656# a_10020_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X7863 VDD buf_in2.inv0.O buf_in2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7864 VSS word8.byte1.tinv3.I a_153300_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7865 word5.byte3.dff_5.O word5.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7866 word4.byte1.dff_6.O word4.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7867 VSS a_144660_5492# word4.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7868 a_147660_4226# a_147430_3276# a_147100_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7869 a_44580_5492# a_44370_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7870 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7871 a_73020_2660# word2.byte3.cgate0.nand0.A word2.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7872 a_47970_3326# a_47350_3276# a_47860_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7873 a_140130_4226# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X7874 buf_in19.inv1.O buf_in19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7875 a_150930_2776# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7876 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7877 a_19380_2356# a_19170_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7878 VDD a_40980_11764# word8.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7879 word2.byte1.dff_6.O word2.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7880 word3.byte3.dff_5.O word3.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7881 VDD a_66180_11764# word8.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X7882 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7883 a_75900_13636# dec8.and4_6.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7884 a_48140_7362# word5.byte3.cgate0.inv1.O a_47970_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7885 word6.byte2.dff_2.O word6.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7886 a_140460_7978# a_140230_8768# a_139900_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7887 VDD word1.byte1.cgate0.nand0.B word1.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7888 a_40770_7978# a_40150_8768# a_40660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7889 word2.byte3.tinv7.O word2.byte3.tinv0.EN a_42420_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7890 a_106680_3442# word3.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7891 VSS word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7892 a_160500_6578# word5.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7893 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7894 VDD word8.byte1.tinv7.I a_167700_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7895 a_144660_10088# a_144450_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7896 word6.byte3.dff_3.O word6.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7897 word1.byte1.tinv7.O buf_out8.inv0.I a_142500_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7898 a_110280_306# word1.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7899 a_48140_4226# word3.byte3.cgate0.inv1.O a_47970_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7900 a_58940_2776# a_58150_2496# a_58770_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7901 word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.latch0.I0.O a_92280_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7902 VDD word1.byte4.tinv5.I a_20820_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7903 a_67620_3442# word3.byte3.tinv7.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7904 VSS a_104080_140# a_103080_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7905 a_111510_9598# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7906 VSS a_48180_6952# word5.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7907 a_15180_190# word1.byte4.cgate0.inv1.O a_14620_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7908 VSS buf_out10.inv0.O buf_out10.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7909 VSS a_106680_4840# a_108240_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7910 a_126520_4842# a_124680_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7911 a_101040_9598# word7.byte2.dff_7.CLK a_100480_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7912 VSS a_48180_3816# word3.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7913 VSS buf_out6.inv0.I buf_out6.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X7914 VSS Di29 buf_in30.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7915 VSS buf_in26.inv0.O buf_in26.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7916 a_25750_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7917 a_51460_2776# a_49620_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7918 a_126520_1706# a_124680_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7919 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7920 a_167700_5796# word4.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7921 VDD buf_out27.inv0.O Do26_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7922 VDD buf_out21.inv0.O Do20_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7923 VDD buf_in8.inv0.O buf_in8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7924 a_155420_11114# word8.byte1.dff_7.CLK a_155250_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7925 a_166220_1090# word1.byte1.dff_7.CLK a_166050_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7926 a_22660_9048# a_20820_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7927 word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.latch0.I0.O a_75720_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7928 word6.gt_re1.O word6.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7929 VSS word1.byte4.inv_and.O a_36120_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7930 word4.byte2.tinv7.O word4.byte2.tinv6.EN a_124680_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7931 a_64020_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7932 VSS a_114880_1656# a_113880_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7933 VSS buf_sel4.inv0.O buf_sel4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7934 VDD word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7935 a_40380_10498# a_40150_9548# a_39820_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7936 VSS a_151860_2356# word2.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7937 a_103080_9714# word7.byte2.tinv0.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7938 VSS word6.byte4.tinv7.I a_28020_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7939 word2.byte4.cgate0.inv1.I word2.byte4.cgate0.nand0.A a_33420_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7940 a_51780_2356# a_51570_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7941 a_128280_7364# word5.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7942 a_4660_1090# a_2820_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7943 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7944 VDD word7.byte1.cgate0.nand0.B word7.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7945 VDD word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7946 a_22980_8628# a_22770_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7947 word5.byte3.inv_and.O word5.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7948 a_19170_4842# a_18550_5632# a_19060_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7949 VSS buf_sel8.inv0.I buf_sel8.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7950 a_162060_11114# a_161830_11904# a_161500_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7951 a_21820_9548# word7.byte4.cgate0.inv1.O a_22050_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X7952 word5.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7953 word1.gt_re3.I word1.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7954 a_128280_4228# word3.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7955 a_122920_11114# a_121080_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X7956 a_154630_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7957 VSS a_143500_9548# a_142500_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X7958 a_55380_6952# a_55170_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7959 VSS word1.byte1.cgate0.nand0.B a_73020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7960 VDD word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7961 a_19170_1706# a_18550_2496# a_19060_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7962 word3.byte3.inv_and.O word3.byte3.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7963 a_166260_6952# a_166050_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7964 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7965 a_18450_2776# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X7966 word3.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7967 VDD a_156900_4840# a_158460_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7968 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7969 a_65350_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7970 VSS word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X7971 a_4980_680# a_4770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7972 a_53220_306# word1.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7973 a_62540_9048# a_61750_8768# a_62370_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X7974 word3.byte4.tinv7.O word3.byte4.tinv7.EN a_28020_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X7975 a_144450_6462# word5.byte1.dff_7.CLK a_144340_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7976 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7977 a_55380_3816# a_55170_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X7978 VDD a_103080_11112# a_104640_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7979 VSS a_112440_10088# word7.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X7980 a_166260_3816# a_166050_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7981 VDD a_156900_1704# a_158460_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7982 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7983 a_65350_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X7984 VDD buf_in9.inv0.O buf_in9.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7985 VDD word6.byte4.nand.OUT word6.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X7986 a_144450_3326# word3.byte1.dff_7.CLK a_144340_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7987 a_105240_5492# a_105030_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X7988 a_115210_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7989 word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.latch0.I0.ENB a_36120_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7990 word7.byte1.inv_and.O word7.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7991 VSS a_113880_1704# a_115440_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7992 VSS buf_in24.inv0.O buf_in24.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7993 VDD a_46020_7976# a_47580_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X7994 a_2820_4840# word4.byte4.tinv0.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X7995 word4.byte4.dff_0.O word4.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X7996 VSS word2.byte1.tinv1.I a_146100_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X7997 VSS a_142500_11112# a_144060_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X7998 VDD buf_in17.inv0.O buf_in17.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X7999 buf_in5.inv0.O Di4 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8000 VSS word8.byte3.tinv2.I a_49620_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8001 VDD word5.byte4.tinv1.I a_6420_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8002 a_55380_680# a_55170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8003 a_105240_2356# a_105030_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8004 a_105030_11114# word8.byte2.dff_7.CLK a_104920_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8005 VSS word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8006 a_33420_306# word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8007 a_126630_4842# word4.byte2.dff_7.CLK a_126520_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8008 a_8370_7978# word6.byte4.cgate0.inv1.O a_8260_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8009 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8010 VDD a_62580_5492# word4.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8011 VSS word8.byte3.cgate0.nand0.A a_75360_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8012 VDD word3.byte4.tinv1.I a_6420_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8013 VDD word5.buf_ck1.I word5.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8014 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8015 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8016 a_10020_11112# word8.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8017 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8018 VDD a_62580_2356# word2.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8019 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.latch0.I0.O a_131700_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8020 a_111280_11064# a_111610_11904# a_111510_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8021 a_22940_190# a_22150_140# a_22770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8022 a_11580_5912# word4.byte4.cgate0.inv1.O a_11020_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8023 VDD word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8024 VDD word3.buf_ck1.I word3.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8025 buf_sel5.inv1.O buf_sel5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8026 VDD word6.byte1.buf_RE1.I word6.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8027 a_49620_6578# buf_out22.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8028 VSS a_4980_2356# a_4940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8029 word8.byte1.dff_6.O word8.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8030 word1.byte4.dff_2.O word1.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8031 a_58380_2776# word2.byte3.cgate0.inv1.O a_57820_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8032 a_111280_6412# a_111610_6412# a_111510_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8033 VDD a_3820_140# a_2820_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8034 word3.byte3.tinv7.O word3.byte3.tinv5.EN a_60420_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8035 a_49620_3442# buf_out22.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8036 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8037 VSS a_144660_11764# word8.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8038 a_11970_9598# word7.byte4.cgate0.inv1.O a_11860_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8039 a_17220_4840# word4.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8040 VSS word8.byte2.tinv3.I a_113880_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8041 a_111280_3276# a_111610_3276# a_111510_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8042 VDD word8.buf_ck1.I word8.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8043 word7.byte4.dff_6.O word7.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8044 a_54450_6462# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8045 VSS buf_in8.inv0.O buf_in8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8046 a_142500_9714# word7.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8047 VSS buf_in29.inv0.O buf_in29.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8048 a_165330_7362# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8049 VDD a_40980_10088# word7.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8050 a_17220_1704# word2.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8051 VSS a_162660_6952# a_162620_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8052 VDD buf_out2.inv0.I buf_out2.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X8053 VDD a_66180_10088# word7.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8054 a_26260_7978# a_24420_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8055 VSS a_25420_140# a_24420_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8056 a_54450_3326# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8057 word2.byte2.buf_RE1.I word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8058 a_4050_7978# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8059 a_12140_9598# a_11350_9548# a_11970_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8060 a_165330_4226# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8061 VDD word8.byte2.tinv7.I a_128280_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8062 VSS buf_ck.inv0.O CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8063 VSS a_162660_3816# a_162620_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8064 a_165660_7978# a_165430_8768# a_165100_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8065 a_105200_5912# a_104410_5632# a_105030_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8066 a_65970_7978# a_65350_8768# a_65860_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8067 a_104310_4842# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8068 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8069 word2.byte3.tinv7.O word2.byte3.tinv7.EN a_67620_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8070 a_14850_12184# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8071 a_151540_9598# a_149700_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8072 VSS word4.byte1.cgate0.nand0.B word4.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8073 VSS a_51780_10088# a_51740_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8074 VDD buf_re.inv1.O word7.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8075 a_26580_8628# a_26370_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8076 word1.byte1.tinv7.O buf_out1.inv0.I a_167700_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8077 VDD word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8078 VDD a_108840_6952# a_108800_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8079 word1.byte1.tinv7.O word1.byte1.tinv4.EN a_156900_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8080 a_58380_11114# a_58150_11904# a_57820_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8081 a_153300_11112# buf_out5.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8082 a_105030_7978# word6.byte2.dff_7.CLK a_104920_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8083 VDD word1.byte2.tinv3.I a_113880_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8084 word7.buf_sel0.O buf_sel7.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X8085 VSS a_14620_4792# a_13620_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8086 VSS a_42420_306# a_43980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8087 a_104310_1706# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8088 word6.byte1.tinv7.O buf_out5.inv0.I a_153300_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8089 a_142500_6578# word5.byte1.tinv0.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8090 buf_sel7.inv1.O buf_sel7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8091 VSS word7.byte3.tinv1.I a_46020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8092 VDD a_108840_3816# a_108800_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8093 VSS word3.byte1.nand.B a_39180_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8094 a_14620_11064# word8.byte4.cgate0.inv1.O a_14850_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8095 a_1340_6462# a_550_6412# a_1170_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8096 a_66140_7978# word6.byte3.cgate0.inv1.O a_65970_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8097 word5.byte4.tinv7.O buf_out30.inv0.I a_10020_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8098 a_92280_6578# word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8099 VSS buf_in9.inv0.O buf_in9.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8100 word7.byte2.tinv7.O buf_out9.inv0.I a_128280_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8101 VDD a_101640_8628# a_101600_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8102 a_1340_3326# a_550_3276# a_1170_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8103 a_58660_12184# a_56820_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8104 word3.byte4.tinv7.O buf_out30.inv0.I a_10020_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8105 a_155420_10498# word7.byte1.dff_7.CLK a_155250_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8106 a_61750_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8107 word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.latch0.I0.O a_93540_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8108 VSS a_3820_1656# a_2820_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8109 VSS buf_out26.inv0.O Do25_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8110 a_95160_8932# word6.byte2.cgate0.nand0.A word6.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8111 word6.byte2.tinv7.O word6.byte2.tinv0.EN a_103080_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8112 word5.byte2.dff_3.O word5.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8113 VDD a_166260_6952# word5.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8114 a_42420_306# word1.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8115 VDD buf_out8.inv0.O Do7_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8116 VDD buf_in20.inv0.O buf_in20.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8117 a_118710_1090# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8118 a_47860_9048# a_46020_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8119 VDD a_44580_11764# a_44540_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8120 a_140230_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8121 VDD a_166260_3816# word3.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8122 word3.byte2.dff_3.O word3.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8123 word4.byte1.dff_2.O word4.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8124 VSS buf_out32.inv0.I buf_out32.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X8125 a_162060_10498# a_161830_9548# a_161500_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8126 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8127 a_115210_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8128 a_122920_10498# a_121080_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8129 a_125680_4792# a_126010_5632# a_125910_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8130 VDD a_105240_5492# word4.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8131 buf_in22.inv1.O buf_in22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8132 a_1340_11114# word8.byte4.cgate0.inv1.O a_1170_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8133 a_140230_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8134 VSS word7.byte1.nand.B a_78780_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8135 VSS word3.byte1.tinv6.I a_164100_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8136 a_48180_8628# a_47970_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8137 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8138 word5.byte1.cgate0.nand0.A word5.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8139 buf_sel1.inv1.O buf_sel1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8140 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8141 a_112400_2776# a_111610_2496# a_112230_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8142 VDD a_49620_11112# a_51180_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8143 VSS a_1380_10088# word7.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8144 VSS a_17220_9714# a_18780_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8145 VDD a_105240_2356# word2.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8146 VDD a_103080_9714# a_104640_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8147 a_131700_4840# word4.byte1.cgate0.latch0.I0.ENB word4.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8148 word5.byte3.cgate0.inv1.I word5.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8149 VSS word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8150 word8.byte3.dff_5.O word8.byte3.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8151 word5.byte2.cgate0.inv1.I word5.byte2.cgate0.nand0.A a_95160_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8152 a_14620_7928# word6.byte4.cgate0.inv1.O a_14850_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8153 a_122410_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8154 a_116000_6462# a_115210_6412# a_115830_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8155 a_131700_1704# word2.byte1.cgate0.latch0.I0.ENB word2.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8156 VSS a_2820_1704# a_4380_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8157 a_550_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8158 word3.byte3.cgate0.inv1.I word3.byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8159 a_64020_7976# word6.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8160 VSS word5.byte3.tinv3.I a_53220_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8161 word4.byte2.cgate0.nand0.A word4.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8162 a_116000_3326# a_115210_3276# a_115830_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8163 a_8580_11764# a_8370_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8164 a_51570_11114# word8.byte3.cgate0.inv1.O a_51460_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8165 a_20820_7976# buf_out27.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8166 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8167 a_11350_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8168 a_128280_306# word1.byte2.tinv7.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8169 word2.byte2.cgate0.nand0.A word2.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8170 VSS buf_in23.inv0.O buf_in23.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8171 buf_re.inv0.O RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8172 a_67620_306# word1.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8173 VDD buf_in4.inv0.O buf_in4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8174 a_10020_11112# word8.byte4.tinv2.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8175 VDD buf_in25.inv0.O buf_in25.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8176 a_151820_1090# word1.byte1.dff_7.CLK a_151650_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8177 VDD a_65020_6412# a_64020_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8178 a_128280_2660# word2.byte2.tinv7.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8179 word4.byte2.tinv7.O word4.byte2.tinv2.EN a_110280_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8180 VSS a_160500_6578# a_162060_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8181 VSS word6.byte4.tinv3.I a_13620_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8182 VDD a_58980_11764# word8.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8183 VSS a_51780_680# a_51740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8184 a_54220_6412# word5.byte3.cgate0.inv1.O a_54450_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8185 a_113880_6578# word5.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8186 VDD a_65020_3276# a_64020_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8187 word2.byte1.dff_4.O word2.byte1.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8188 VSS a_160500_3442# a_162060_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8189 VSS word8.byte3.buf_RE0.O word8.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8190 word8.byte2.dff_6.O word8.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8191 buf_sel7.inv1.O buf_sel7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8192 a_108630_7978# a_108010_8768# a_108520_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8193 a_18550_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8194 a_113880_3442# word3.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8195 a_54220_3276# word3.byte3.cgate0.inv1.O a_54450_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8196 VSS a_49620_9714# a_51180_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8197 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8198 word4.byte4.dff_4.O word4.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8199 a_104080_7928# a_104410_8768# a_104310_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8200 VSS a_105240_11764# word8.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8201 VSS word7.buf_ck1.I word7.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8202 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8203 a_50950_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8204 a_103080_9714# word7.byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8205 word2.byte4.dff_4.O word2.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8206 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8207 VSS buf_in16.inv0.O buf_in16.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8208 VDD word1.byte4.nand.OUT word1.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8209 VDD word4.byte3.dff_0.O_bar a_42420_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8210 a_26260_11114# a_24420_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8211 word6.gt_re3.I word6.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8212 a_4980_680# a_4770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8213 a_148220_6462# a_147430_6412# a_148050_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8214 a_47250_9048# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8215 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8216 word7.byte2.dff_4.O word7.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8217 a_13620_6578# word5.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8218 a_50950_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8219 VDD buf_out10.inv0.I buf_out10.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X8220 VDD word8.gt_re1.O word8.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8221 a_100810_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8222 VSS word1.byte1.nand.B a_78780_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8223 VSS buf_out8.inv0.I buf_out8.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X8224 VSS a_155460_8628# a_155420_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8225 VSS a_105240_680# word1.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8226 VDD word2.byte3.dff_0.O_bar a_42420_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8227 VSS buf_in28.inv0.O buf_in28.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8228 VSS buf_out1.inv0.I buf_out1.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X8229 a_148220_3326# a_147430_3276# a_148050_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8230 a_144340_4842# a_142500_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8231 VDD a_44580_5492# a_44540_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8232 VSS word2.byte1.inv_and.O a_131700_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8233 a_119320_2776# a_117480_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8234 VDD buf_out23.inv0.O Do22_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8235 VDD buf_in3.inv0.O buf_in3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8236 a_144340_1706# a_142500_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8237 word1.byte3.dff_0.O word1.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8238 VDD a_44580_2356# a_44540_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8239 buf_in22.inv1.O buf_in22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8240 VDD word7.byte3.dff_0.O_bar a_42420_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8241 VSS word4.byte1.cgate0.nand0.B word4.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8242 a_58380_10498# a_58150_9548# a_57820_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8243 word2.byte2.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B a_93540_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8244 word6.byte4.dff_1.O word6.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8245 a_2820_3442# word3.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8246 word4.byte1.tinv7.O word4.byte1.tinv0.EN a_142500_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8247 dec8.and4_0.nand1.OUT dec8.and4_3.nand1.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8248 VSS a_48180_5492# word4.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8249 VSS a_65020_7928# a_64020_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8250 word7.byte2.tinv7.O word7.byte2.tinv5.EN a_121080_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8251 a_39180_2660# buf_we1.inv1.O word2.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8252 VSS word4.byte4.tinv5.I a_20820_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8253 a_154860_11114# a_154630_11904# a_154300_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8254 a_14620_9548# word7.byte4.cgate0.inv1.O a_14850_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8255 VDD word1.byte1.buf_RE1.I word1.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8256 a_146100_6578# word5.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8257 a_73560_12850# dec8.and4_5.nand1.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8258 a_119040_4842# a_118810_5632# a_118480_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8259 word6.byte1.dff_5.O word6.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8260 a_39180_306# buf_we1.inv1.O word1.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8261 a_167700_6578# word5.byte1.tinv7.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8262 a_19340_1090# word1.byte4.cgate0.inv1.O a_19170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8263 VDD word6.byte2.tinv6.I a_124680_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8264 buf_sel8.inv1.O buf_sel8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8265 word8.byte4.dff_7.O word8.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8266 VSS word7.gt_re1.O word7.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8267 a_146100_3442# word3.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8268 VSS word3.byte3.inv_and.O a_75720_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8269 VDD word5.byte4.cgate0.nand0.A a_35760_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8270 a_43980_2776# word2.byte3.cgate0.inv1.O a_43420_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8271 a_119040_1706# a_118810_2496# a_118480_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8272 a_154300_140# a_154630_140# a_154530_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8273 a_7750_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8274 a_26580_11764# a_26370_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8275 a_61750_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8276 a_158740_1090# a_156900_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8277 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8278 a_75720_6578# word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8279 VDD a_58980_680# a_58940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8280 VDD a_126840_8628# a_126800_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8281 VDD a_14620_9548# a_13620_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8282 VSS word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8283 VDD word3.byte4.cgate0.nand0.A a_35760_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8284 VDD a_125680_7928# a_124680_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8285 VDD a_21820_4792# a_20820_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8286 VDD buf_out16.inv0.O buf_out16.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8287 word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.latch0.I0.O a_75720_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8288 VDD a_44580_10088# a_44540_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8289 a_10020_1704# word2.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8290 VSS buf_out7.inv0.O Do6_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8291 word6.byte2.tinv7.O word6.byte2.tinv7.EN a_128280_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8292 VDD a_21820_1656# a_20820_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8293 a_150930_7362# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8294 a_19380_6952# a_19170_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8295 a_1340_10498# word7.byte4.cgate0.inv1.O a_1170_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8296 a_11860_7978# a_10020_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8297 a_22150_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8298 VDD a_166260_11764# a_166220_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8299 a_57820_9548# a_58150_9548# a_58050_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8300 a_78780_8932# buf_we2.inv1.O word6.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8301 VSS word6.byte2.nand.OUT word6.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8302 a_55380_5492# a_55170_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8303 a_165430_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8304 a_164100_1704# word2.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8305 a_150930_4226# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8306 a_151260_1090# a_151030_140# a_150700_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8307 a_19380_3816# a_19170_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8308 a_51570_190# a_50950_140# a_51460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8309 VDD a_49620_9714# a_51180_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8310 a_36120_8932# word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8311 a_58940_7362# word5.byte3.cgate0.inv1.O a_58770_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8312 a_22150_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8313 word4.gt_re3.I word4.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8314 Do21_buf buf_out22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8315 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8316 a_165430_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8317 a_162620_4842# word4.byte1.dff_7.CLK a_162450_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8318 a_144450_4842# word4.byte1.dff_7.CLK a_144340_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8319 word1.byte3.dff_6.O word1.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8320 word2.byte3.tinv7.O word2.byte3.tinv3.EN a_53220_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8321 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8322 a_12180_8628# a_11970_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8323 word1.byte1.tinv7.O buf_out5.inv0.I a_153300_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8324 VDD word8.byte1.cgate0.nand0.B word8.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8325 a_155460_10088# a_155250_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8326 a_126240_190# word1.byte2.dff_7.CLK a_125680_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8327 VSS a_55380_2356# word2.byte3.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8328 a_58940_4226# word3.byte3.cgate0.inv1.O a_58770_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8329 a_54550_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8330 a_162620_1706# word2.byte1.dff_7.CLK a_162450_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8331 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8332 a_156900_4840# buf_out4.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8333 a_53220_4840# word4.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8334 a_107680_7928# word6.byte2.dff_7.CLK a_107910_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8335 VDD word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8336 a_108800_9048# a_108010_8768# a_108630_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8337 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8338 VSS a_26580_8628# word6.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8339 a_8580_10088# a_8370_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8340 a_160500_11112# word8.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8341 a_51740_7978# word6.byte3.cgate0.inv1.O a_51570_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8342 VDD word6.byte1.tinv4.I a_156900_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8343 VSS a_58980_6952# word5.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8344 a_156900_1704# buf_out4.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8345 a_36120_3442# word3.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8346 VDD word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8347 word5.byte2.inv_and.O word5.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8348 word6.byte4.cgate0.nand0.A word6.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8349 a_51460_7362# a_49620_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8350 VDD a_8580_680# word1.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8351 VDD buf_in12.inv0.O buf_in12.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8352 VSS word8.byte2.tinv1.I a_106680_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8353 word4.byte3.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8354 a_46020_7976# buf_out23.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8355 word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.latch0.I0.O a_36120_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8356 VSS a_58980_3816# word3.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8357 a_1380_5492# a_1170_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8358 a_104410_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8359 VDD a_159060_8628# a_159020_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8360 VDD word8.byte2.buf_RE1.I word8.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8361 a_51460_4226# a_49620_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8362 VSS buf_in3.inv0.O buf_in3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8363 word7.byte4.tinv7.O buf_out26.inv0.I a_24420_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8364 word2.byte3.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8365 VDD a_151860_6952# word5.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8366 VDD a_58980_10088# word7.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8367 a_160500_7976# word6.byte1.tinv5.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8368 a_1380_2356# a_1170_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8369 VDD buf_in8.inv0.O buf_in8.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8370 a_131700_12068# word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8371 a_51780_6952# a_51570_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8372 VSS word8.byte4.nand.OUT word8.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8373 VDD a_42420_4840# a_43980_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8374 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8375 buf_we2.inv1.O buf_we2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8376 VDD a_151860_3816# word3.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8377 a_18550_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8378 word6.byte4.dff_2.O word6.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8379 VSS a_12180_2356# a_12140_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8380 a_51780_3816# a_51570_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8381 VDD a_42420_1704# a_43980_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8382 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8383 buf_in18.inv1.O buf_in18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8384 a_111280_4792# a_111610_5632# a_111510_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8385 VSS word8.byte4.buf_RE0.O word8.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8386 a_101640_8628# a_101430_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8387 VSS a_220_140# a_120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8388 VDD a_11020_140# a_10020_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8389 VSS word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8390 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8391 buf_sel8.inv1.O buf_sel8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8392 a_146100_11112# buf_out7.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8393 a_18450_7362# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8394 VSS a_26580_680# word1.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8395 a_144340_190# a_142500_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8396 a_151650_1706# word2.byte1.dff_7.CLK a_151540_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8397 VSS a_15780_6952# a_15740_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8398 a_149700_3442# word3.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8399 a_54450_5912# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8400 VSS word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8401 a_26260_10498# a_24420_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8402 word3.byte2.tinv7.O word3.byte2.tinv1.EN a_106680_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8403 VSS word3.byte2.buf_RE1.I word3.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8404 a_18450_4226# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8405 word7.byte2.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8406 a_64020_306# word1.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8407 VSS a_15780_3816# a_15740_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8408 VSS a_162660_5492# a_162620_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8409 word5.byte1.tinv7.O word5.byte1.tinv5.EN a_160500_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8410 VSS buf_out16.inv0.I buf_out16.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X8411 a_18780_7978# a_18550_8768# a_18220_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8412 VDD word4.byte3.tinv7.I a_67620_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8413 VDD a_113880_6578# a_115440_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8414 a_20820_306# buf_out27.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8415 a_43650_11114# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8416 a_11250_7978# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8417 a_8260_2776# a_6420_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8418 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8419 a_154530_9598# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8420 VSS a_111280_140# a_110280_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8421 a_108800_11114# word8.byte2.dff_7.CLK a_108630_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8422 VDD a_56820_306# a_58380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8423 VSS word1.byte1.buf_RE0.I word1.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8424 word8.byte3.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8425 VDD word2.byte3.tinv7.I a_67620_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8426 VDD a_113880_3442# a_115440_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8427 a_112230_9598# word7.byte2.dff_7.CLK a_112120_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8428 a_22380_190# word1.byte4.cgate0.inv1.O a_21820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8429 VSS a_1380_680# a_1340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8430 word5.byte4.dff_5.O word5.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8431 a_8580_2356# a_8370_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8432 VDD a_50620_6412# a_49620_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8433 a_113880_1704# word2.byte2.tinv3.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8434 VDD word7.byte1.tinv6.I a_164100_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8435 a_7980_4842# a_7750_5632# a_7420_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8436 dec8.and4_2.nand1.OUT dec8.and4_3.nand1.A a_68160_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8437 buf_in2.inv1.O buf_in2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8438 a_154860_10498# a_154630_9548# a_154300_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8439 word3.byte4.dff_5.O word3.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8440 a_1340_5912# a_550_5632# a_1170_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8441 word4.byte1.tinv7.O word4.byte1.tinv7.EN a_167700_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8442 VSS word4.byte2.tinv3.I a_113880_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8443 a_42420_11112# word8.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8444 VDD a_50620_3276# a_49620_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8445 VDD buf_in31.inv0.O buf_in31.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8446 buf_in17.inv1.O buf_in17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8447 word7.byte4.dff_7.O word7.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8448 a_146100_9714# word7.byte1.tinv1.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8449 VDD a_4980_6952# a_4940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8450 a_75720_2660# word2.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8451 a_7980_1706# a_7750_2496# a_7420_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8452 a_58380_7362# a_58150_6412# a_57820_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8453 a_162060_4842# a_161830_5632# a_161500_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8454 a_62370_4842# a_61750_5632# a_62260_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8455 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8456 VSS word2.byte1.cgate0.nand0.B a_33420_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8457 VDD a_4980_3816# a_4940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8458 a_75360_12068# word8.byte1.cgate0.nand0.B word8.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8459 word8.byte1.dff_2.O word8.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8460 a_162060_1706# a_161830_2496# a_161500_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8461 VSS a_11020_1656# a_10020_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8462 a_58380_4226# a_58150_3276# a_57820_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8463 a_55060_9598# a_53220_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8464 a_62370_1706# a_61750_2496# a_62260_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8465 word4.byte1.tinv7.O buf_out6.inv0.I a_149700_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8466 VDD word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8467 a_56820_11112# word8.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8468 word1.gt_re3.I word1.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8469 a_61650_2776# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8470 VSS word1.byte1.tinv0.I a_142500_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8471 VSS word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8472 a_51180_7978# a_50950_8768# a_50620_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8473 a_140230_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8474 word2.byte1.tinv7.O buf_out6.inv0.I a_149700_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8475 VDD word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8476 VSS word3.byte4.tinv4.I a_17220_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8477 a_28020_4840# word4.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8478 buf_in15.inv0.O buf_in15.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8479 word7.byte2.dff_0.O word7.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8480 VSS a_155460_10088# word7.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8481 word6.byte3.tinv7.O word6.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8482 VSS word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8483 VDD a_101640_11764# a_101600_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8484 VDD a_166260_10088# a_166220_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8485 a_47580_190# word1.byte3.cgate0.inv1.O a_47020_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8486 VSS buf_out29.inv0.O Do28_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8487 buf_in6.inv0.O Di5 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8488 VSS a_220_7928# a_120_7978# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8489 a_122640_6462# word5.byte2.dff_7.CLK a_122080_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8490 a_158230_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8491 a_28020_1704# word2.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8492 a_148260_5492# a_148050_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8493 VDD buf_re.inv0.O buf_re.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8494 a_28020_12068# word8.byte4.tinv7.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8495 a_104920_2776# a_103080_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8496 a_47350_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8497 a_22940_9598# a_22150_9548# a_22770_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8498 a_122640_3326# word3.byte2.dff_7.CLK a_122080_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8499 VDD word8.byte1.nand.B word8.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8500 a_148260_2356# a_148050_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8501 Do20_buf buf_out21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8502 VSS word6.byte1.cgate0.nand0.B a_73020_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8503 a_47350_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8504 a_116000_5912# a_115210_5632# a_115830_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8505 VSS a_6420_11112# a_7980_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8506 VSS a_50620_7928# a_49620_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8507 a_6420_6578# buf_out31.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8508 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8509 VSS word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8510 a_131700_7364# word5.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8511 VDD word1.byte2.tinv6.I a_124680_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8512 a_121080_11112# word8.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8513 word3.byte1.inv_and.O word3.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8514 a_6420_3442# buf_out31.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8515 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8516 VDD word5.buf_ck1.I word5.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8517 a_150700_1656# a_151030_2496# a_150930_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8518 buf_sel7.inv1.O buf_sel7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8519 VSS word7.byte3.tinv4.I a_56820_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8520 VSS a_117480_9714# a_119040_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8521 VSS a_13620_6578# a_15180_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8522 a_131700_4228# word3.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8523 VSS a_165100_6412# a_164100_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8524 a_93540_7364# word5.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8525 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8526 VSS word1.byte1.tinv7.I a_167700_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8527 word8.byte4.cgate0.nand0.A word8.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8528 VDD a_112440_680# a_112400_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8529 VDD word3.buf_ck1.I word3.byte1.cgate0.nand0.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8530 VSS buf_in11.inv0.O buf_in11.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8531 VSS a_13620_3442# a_15180_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8532 VSS a_160500_4840# a_162060_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8533 a_11020_4792# word4.byte4.cgate0.inv1.O a_11250_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8534 a_154300_6412# a_154630_6412# a_154530_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8535 VSS a_165100_3276# a_164100_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8536 VDD buf_out12.inv0.I buf_out12.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X8537 a_93540_4228# word3.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8538 a_73020_6578# word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8539 a_60420_4840# word4.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8540 VDD word8.byte3.tinv5.I a_60420_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8541 a_11020_1656# word2.byte4.cgate0.inv1.O a_11250_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8542 VDD word6.byte4.buf_RE0.O word6.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8543 a_154300_3276# a_154630_3276# a_154530_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8544 VSS a_54220_9548# a_53220_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8545 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8546 a_60420_1704# word2.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8547 VDD buf_in28.inv0.O buf_in28.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8548 a_43420_9548# a_43750_9548# a_43650_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8549 VSS word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8550 VSS buf_in31.inv0.O buf_in31.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8551 VSS Di4 buf_in5.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8552 a_6420_9714# word7.byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8553 buf_in17.inv1.O buf_in17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8554 a_106680_11112# buf_out15.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8555 VSS a_8580_10088# a_8540_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8556 a_112400_7362# word5.byte2.dff_7.CLK a_112230_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8557 buf_in22.inv1.O buf_in22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8558 VSS word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8559 a_126840_8628# a_126630_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8560 VDD a_116040_5492# word4.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8561 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8562 a_780_6462# word5.byte4.cgate0.inv1.O a_220_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8563 a_112400_4226# word3.byte2.dff_7.CLK a_112230_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8564 a_148220_5912# a_147430_5632# a_148050_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8565 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8566 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8567 a_147330_4842# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8568 VSS buf_out20.inv0.O Do19_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8569 VDD a_2820_6578# a_4380_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8570 a_119430_190# word1.byte2.dff_7.CLK a_119320_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8571 VSS a_40980_2356# word2.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8572 VDD a_116040_2356# word2.byte2.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8573 a_25420_140# word1.byte4.cgate0.inv1.O a_25650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8574 VSS word8.byte2.buf_RE1.I word8.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8575 VDD word5.gt_re1.O word5.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8576 VDD word1.byte1.tinv4.I a_156900_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8577 buf_sel6.inv0.I dec8.and4_5.nand1.OUT a_74100_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8578 a_43650_10498# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8579 a_148050_7978# word6.byte1.dff_7.CLK a_147940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8580 a_780_3326# word3.byte4.cgate0.inv1.O a_220_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8581 word7.byte1.tinv7.O word7.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8582 a_147330_1706# buf_in6.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8583 VSS word4.byte4.nand.OUT word4.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8584 a_108800_10498# word7.byte2.dff_7.CLK a_108630_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8585 VDD word5.byte4.buf_RE0.O word5.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8586 word1.byte4.cgate0.nand0.A word1.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8587 word1.byte1.tinv7.O word1.byte1.tinv6.EN a_164100_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8588 VDD a_2820_3442# a_4380_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8589 a_19380_11764# a_19170_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8590 a_1170_9598# word7.byte4.cgate0.inv1.O a_1060_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8591 VDD word6.byte1.tinv0.I a_142500_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8592 VSS word7.buf_sel0.O word7.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8593 VSS word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8594 VDD word3.gt_re1.O word3.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8595 a_46020_306# buf_out23.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8596 VSS a_49620_306# a_51180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8597 a_11970_11114# a_11350_11904# a_11860_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8598 a_165940_12184# a_164100_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8599 a_165330_11114# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8600 VDD word6.byte2.inv_and.O a_92280_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8601 VDD word3.byte4.buf_RE0.O word3.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8602 VDD a_144660_8628# a_144620_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8603 word6.byte4.dff_3.O word6.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8604 a_151030_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8605 VSS word6.byte1.cgate0.nand0.B a_134580_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8606 word5.byte3.dff_1.O word5.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8607 VSS a_139800_7978# a_140460_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8608 VDD buf_out25.inv0.O Do24_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8609 word5.byte1.dff_4.O word5.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8610 word6.byte1.tinv7.O word6.byte1.tinv1.EN a_146100_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8611 a_110280_306# word1.byte2.tinv2.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8612 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8613 buf_in23.inv1.O buf_in23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8614 word3.byte3.dff_1.O word3.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8615 a_22380_9598# word7.byte4.cgate0.inv1.O a_21820_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8616 VSS word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8617 word3.byte1.dff_4.O word3.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8618 VSS word4.byte1.buf_RE1.I word4.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8619 VDD buf_out31.inv0.O Do30_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8620 VSS a_57820_140# a_56820_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8621 a_164100_11112# word8.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8622 a_119430_190# a_118810_140# a_119320_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8623 word7.byte1.dff_2.O word7.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8624 VDD a_148260_5492# word4.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8625 VDD word8.byte4.tinv4.I a_17220_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8626 VDD a_164100_11112# a_165660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8627 a_155420_2776# a_154630_2496# a_155250_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8628 buf_sel3.inv1.O buf_sel3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8629 a_18550_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8630 a_17220_1704# word2.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8631 VSS CLK word7.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8632 VDD a_148260_2356# word2.byte1.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8633 a_134580_6578# word5.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8634 VDD word7.byte1.nand.B word7.byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8635 VDD a_101640_10088# a_101600_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8636 VDD word4.byte2.tinv5.I a_121080_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8637 word8.byte3.tinv7.O buf_out24.inv0.I a_42420_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8638 buf_in14.inv0.O buf_in14.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8639 a_15740_4842# word4.byte4.cgate0.inv1.O a_15570_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8640 VSS word5.gt_re1.O word5.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8641 a_18550_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8642 a_165430_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8643 a_58050_9048# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8644 a_159020_6462# a_158230_6412# a_158850_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8645 word7.byte2.dff_7.O word7.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8646 VDD word2.byte2.tinv5.I a_121080_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8647 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8648 a_119320_7362# a_117480_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8649 a_115440_9048# word6.byte2.dff_7.CLK a_114880_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8650 VDD a_123240_5492# a_123200_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8651 a_15740_1706# word2.byte4.cgate0.inv1.O a_15570_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8652 a_75720_11112# word8.byte3.cgate0.latch0.I0.ENB word8.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8653 word7.byte4.tinv7.O buf_out28.inv0.I a_17220_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8654 a_159020_3326# a_158230_3276# a_158850_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8655 VDD a_122080_4792# a_121080_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8656 word6.byte3.tinv7.O buf_out18.inv0.I a_64020_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8657 a_53220_6578# word5.byte3.tinv3.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8658 a_15570_190# word1.byte4.cgate0.inv1.O a_15460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8659 a_119320_4226# a_117480_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8660 VDD a_123240_2356# a_123200_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8661 VDD buf_in3.inv0.O buf_in3.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8662 VSS word1.byte1.cgate0.inv1.I word1.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8663 VDD a_122080_1656# a_121080_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8664 word1.byte2.dff_2.O word1.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8665 a_112120_7978# a_110280_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8666 word4.byte1.tinv7.O word4.byte1.tinv3.EN a_153300_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8667 VDD Di0 buf_in1.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8668 VSS a_6420_9714# a_7980_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8669 VSS a_58980_5492# word4.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8670 VSS a_44580_11764# word8.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8671 a_56820_7976# word6.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8672 a_75720_10500# word7.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8673 a_43980_7362# a_43750_6412# a_43420_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8674 a_156900_6578# word5.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8675 word8.byte4.tinv7.O word8.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8676 a_3820_7928# word6.byte4.cgate0.inv1.O a_4050_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8677 a_13620_7976# word6.byte4.tinv3.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8678 a_7750_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8679 a_4940_9048# a_4150_8768# a_4770_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8680 word5.byte2.tinv7.O buf_out13.inv0.I a_113880_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8681 a_151860_6952# a_151650_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8682 VDD dec8.and4_5.nand1.B dec8.and4_0.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8683 VDD a_15780_8628# word6.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8684 a_156900_3442# word3.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8685 a_43980_4226# a_43750_3276# a_43420_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8686 a_40660_9598# a_39720_9598# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8687 a_7750_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8688 a_147100_7928# a_147430_8768# a_147330_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8689 a_151860_3816# a_151650_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8690 word3.byte2.tinv7.O buf_out13.inv0.I a_113880_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8691 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8692 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8693 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8694 buf_sel5.inv0.O buf_sel5.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8695 VDD buf_in15.inv0.O buf_in15.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8696 VSS a_141060_10088# word7.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8697 a_550_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8698 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8699 word6.byte1.cgate0.inv1.I word6.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8700 word5.byte4.cgate0.inv1.I word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8701 VDD word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8702 a_40980_10088# a_40770_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8703 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8704 VSS buf_in13.inv0.I buf_in13.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8705 a_42420_4840# buf_out24.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8706 VSS buf_in27.inv0.O buf_in27.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8707 a_22660_1090# a_20820_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8708 a_143830_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8709 VDD a_142500_7976# a_144060_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8710 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8711 VDD a_4980_5492# word4.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8712 VDD word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8713 word3.byte4.cgate0.inv1.I word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8714 word5.byte4.tinv7.O word5.byte4.tinv3.EN a_13620_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8715 VSS a_15780_5492# a_15740_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8716 a_101040_11114# a_100810_11904# a_100480_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8717 a_42420_1704# buf_out24.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8718 a_20820_9714# buf_out27.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8719 VSS a_112440_680# word1.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8720 a_126240_11114# a_126010_11904# a_125680_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8721 VDD a_118480_6412# a_117480_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8722 VDD a_4980_2356# word2.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8723 word1.byte2.tinv7.O word1.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8724 VDD a_55380_6952# word5.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8725 a_131700_2660# word2.byte1.cgate0.latch0.I0.O word2.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8726 a_22980_680# a_22770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8727 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8728 VDD a_118480_3276# a_117480_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8729 buf_in19.inv0.O Di18 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8730 VDD a_55380_3816# word3.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8731 a_140460_12184# word8.byte1.dff_7.CLK a_139900_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8732 word7.byte1.tinv7.O word7.byte1.tinv6.EN a_164100_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8733 word1.byte4.tinv7.O word1.byte4.tinv4.EN a_17220_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8734 a_66140_190# a_65350_140# a_65970_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8735 word2.byte2.cgate0.nand0.A word2.byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8736 VSS word7.byte2.tinv2.I a_110280_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8737 a_64020_4840# word4.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8738 a_100710_11114# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8739 a_118480_7928# word6.byte2.dff_7.CLK a_118710_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8740 word3.byte4.tinv7.O word3.byte4.tinv0.EN a_2820_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8741 dec8.and4_7.nand0.OUT A0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8742 a_11970_9598# a_11350_9548# a_11860_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8743 a_62540_1090# word1.byte3.cgate0.inv1.O a_62370_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8744 a_126520_12184# a_124680_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8745 VSS a_103080_9714# a_104640_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8746 a_165330_10498# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8747 a_20820_4840# word4.byte4.tinv5.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8748 VSS a_150700_6412# a_149700_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8749 word8.byte4.dff_3.O word8.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8750 VDD word7.buf_ck1.I word7.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8751 VDD word6.byte1.tinv7.I a_167700_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8752 word4.byte4.dff_5.O word4.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8753 a_19060_6462# a_17220_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8754 a_55170_1706# word2.byte3.cgate0.inv1.O a_55060_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8755 VSS word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8756 a_124680_7976# buf_out10.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8757 VDD word5.byte4.tinv6.I a_24420_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8758 a_115210_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8759 word2.byte3.dff_7.O word2.byte3.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8760 VSS a_150700_3276# a_149700_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8761 VSS a_106680_11112# a_108240_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8762 a_26370_7978# word6.byte4.cgate0.inv1.O a_26260_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8763 VSS word3.byte1.cgate0.nand0.B word3.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8764 VSS a_119640_6952# word5.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8765 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8766 VDD word1.byte4.buf_RE0.O word1.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8767 a_19060_3326# a_17220_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8768 VDD word4.byte4.cgate0.nand0.A word4.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8769 a_15180_4842# a_14950_5632# a_14620_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8770 VDD a_119640_11764# a_119600_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8771 a_75360_7976# word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8772 a_161500_140# a_161830_140# a_161730_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8773 a_158460_6462# word5.byte1.dff_7.CLK a_157900_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8774 a_58770_6462# word5.byte3.cgate0.inv1.O a_58660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8775 VDD word3.byte4.tinv6.I a_24420_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8776 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8777 VDD word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8778 VSS a_164100_7976# a_165660_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8779 VDD a_12180_6952# a_12140_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8780 VSS a_119640_3816# word3.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8781 a_8370_190# a_7750_140# a_8260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8782 VDD word2.byte4.cgate0.nand0.A word2.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8783 a_15180_1706# a_14950_2496# a_14620_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8784 a_151860_11764# a_151650_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8785 a_158460_3326# word3.byte1.dff_7.CLK a_157900_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8786 VDD buf_out6.inv0.O Do5_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8787 a_58770_3326# word3.byte3.cgate0.inv1.O a_58660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8788 VDD a_53220_4840# a_54780_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8789 VSS word6.byte2.tinv4.I a_117480_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8790 a_61420_11064# a_61750_11904# a_61650_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8791 buf_in5.inv1.O buf_in5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8792 VDD a_12180_3816# a_12140_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8793 word6.byte1.nand.OUT buf_we4.inv1.O a_129540_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8794 VSS a_22980_2356# a_22940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8795 a_151650_6462# a_151030_6412# a_151540_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8796 a_47580_9598# word7.byte3.cgate0.inv1.O a_47020_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8797 VDD a_164100_9714# a_165660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8798 VDD a_12180_11764# word8.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8799 VDD a_53220_1704# a_54780_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8800 buf_in26.inv1.O buf_in26.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8801 buf_in8.inv1.O buf_in8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8802 a_112440_8628# a_112230_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8803 VDD a_4980_11764# a_4940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8804 word8.byte4.inv_and.O word8.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8805 word6.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8806 VDD a_21820_140# a_20820_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8807 VSS a_66180_8628# a_66140_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8808 VSS word6.byte1.cgate0.nand0.B word6.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8809 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8810 a_4940_190# a_4150_140# a_4770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8811 a_151650_3326# a_151030_3276# a_151540_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8812 a_113880_11112# word8.byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8813 VSS a_118480_7928# a_117480_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8814 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8815 a_8540_7978# word6.byte4.cgate0.inv1.O a_8370_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8816 VSS word6.byte4.inv_and.O a_36120_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8817 VSS word2.byte3.dff_0.O_bar a_42420_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8818 word4.gt_re3.I word4.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8819 buf_sel4.inv1.O buf_sel4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8820 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8821 VDD word1.byte1.tinv0.I a_142500_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8822 a_107910_2776# buf_in14.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8823 VSS word8.byte3.tinv6.I a_64020_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8824 a_8260_7362# a_6420_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8825 a_4380_9048# word6.byte4.cgate0.inv1.O a_3820_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8826 a_122640_5912# word4.byte2.dff_7.CLK a_122080_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8827 VSS buf_sel8.inv0.O buf_sel8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8828 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8829 VDD word1.byte2.inv_and.O a_92280_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8830 a_42420_306# word1.byte3.tinv0.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8831 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8832 a_117480_6578# word5.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8833 a_8260_4226# a_6420_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8834 VDD buf_ck.inv0.O CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8835 a_22050_7978# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8836 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8837 a_129540_6578# word5.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8838 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8839 a_8580_6952# a_8370_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8840 VDD word7.byte1.buf_RE1.I word7.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8841 a_123030_9598# word7.byte2.dff_7.CLK a_122920_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8842 word3.byte4.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8843 a_1060_7978# a_120_7978# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8844 VDD a_126840_11764# word8.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8845 a_147430_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8846 VSS a_7420_140# a_6420_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8847 VSS a_18220_6412# a_17220_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8848 a_8580_3816# a_8370_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8849 VDD buf_in9.inv0.I buf_in9.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8850 VDD word7.byte1.cgate0.nand0.B word7.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8851 VSS a_13620_4840# a_15180_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8852 Do23_buf buf_out24.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8853 VDD word7.byte4.inv_and.O a_36120_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8854 VSS a_18220_3276# a_17220_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8855 VSS word4.byte2.tinv6.I a_124680_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8856 Do4_buf buf_out5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8857 a_105030_190# a_104410_140# a_104920_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8858 buf_in17.inv1.O buf_in17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8859 VSS a_139900_1656# a_139800_1706# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8860 a_154300_4792# a_154630_5632# a_154530_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8861 VSS buf_out22.inv0.O Do21_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8862 a_144660_8628# a_144450_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8863 a_68160_12850# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8864 a_61650_7362# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8865 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8866 a_141020_2776# a_140230_2496# a_140850_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8867 VSS a_108840_2356# word2.byte2.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8868 a_40940_11114# word8.byte3.cgate0.inv1.O a_40770_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8869 VSS a_21820_1656# a_20820_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8870 a_66140_11114# word8.byte3.cgate0.inv1.O a_65970_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8871 a_65860_9598# a_64020_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8872 VSS a_125680_4792# a_124680_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8873 a_149700_3442# word3.byte1.tinv2.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8874 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8875 VDD word5.buf_sel0.O word5.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8876 a_61650_4226# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8877 a_151540_190# a_149700_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8878 a_67620_306# word1.byte3.tinv7.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8879 a_18220_11064# a_18550_11904# a_18450_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8880 a_111510_9048# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8881 a_106680_4840# word4.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8882 VDD word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8883 a_61980_7978# a_61750_8768# a_61420_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8884 a_160500_7976# word6.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8885 VSS word7.byte4.cgate0.latch0.I0.O word7.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8886 VDD word3.buf_sel0.O word3.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8887 VSS word5.byte3.buf_RE0.O word5.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8888 a_104920_7362# a_103080_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8889 a_82020_6578# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8890 word1.byte3.tinv7.O buf_out18.inv0.I a_64020_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8891 a_66180_10088# a_65970_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8892 a_101040_9048# word6.byte2.dff_7.CLK a_100480_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8893 a_106680_1704# word2.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8894 VDD word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8895 a_101040_10498# a_100810_9548# a_100480_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8896 VDD word7.byte2.tinv4.I a_117480_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8897 VDD a_7420_6412# a_6420_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8898 buf_in12.inv1.O buf_in12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8899 a_126240_10498# a_126010_9548# a_125680_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8900 a_47860_1090# a_46020_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8901 a_67620_4840# buf_out17.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8902 a_65350_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8903 a_126010_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8904 a_780_5912# word4.byte4.cgate0.inv1.O a_220_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8905 a_104920_4226# a_103080_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X8906 a_101600_9598# a_100810_9548# a_101430_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8907 a_155250_9598# word7.byte1.dff_7.CLK a_155140_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8908 a_48180_11764# a_47970_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8909 VSS a_19380_10088# word7.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8910 VDD a_7420_3276# a_6420_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8911 a_67620_1704# buf_out17.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8912 VSS a_22980_11764# a_22940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8913 a_142500_9714# buf_out8.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X8914 a_126010_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X8915 Do28_buf buf_out29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8916 VSS a_48180_11764# a_48140_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8917 a_39820_6412# a_40150_6412# a_40050_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8918 a_156900_1704# word2.byte1.tinv4.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8919 a_110280_7976# word6.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8920 a_48180_680# a_47970_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8921 buf_in1.inv1.O buf_in1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8922 a_156900_11112# word8.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8923 a_116040_8628# a_115830_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8924 word8.byte4.tinv7.O word8.byte4.tinv5.EN a_20820_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8925 a_100710_10498# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X8926 VSS a_20820_1704# a_22380_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8927 buf_in23.inv1.O buf_in23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8928 a_150700_6412# word5.byte1.dff_7.CLK a_150930_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8929 VDD word7.byte4.dff_0.O_bar a_2820_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8930 VSS word4.byte1.tinv4.I a_156900_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8931 a_39820_3276# a_40150_3276# a_40050_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8932 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8933 word4.byte4.cgate0.nand0.A word4.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8934 a_148260_680# a_148050_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X8935 a_150700_3276# word3.byte1.dff_7.CLK a_150930_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8936 a_161500_1656# a_161830_2496# a_161730_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8937 word2.byte3.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8938 a_46020_4840# word4.byte3.tinv1.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8939 VDD word7.gt_re0.OUT word7.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8940 word4.byte3.dff_1.O word4.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8941 buf_ck.inv0.O buf_ck.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8942 VDD word8.byte4.cgate0.nand0.A a_35760_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8943 VSS a_58980_680# word1.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8944 VDD a_119640_10088# a_119600_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8945 VSS a_112440_8628# word6.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8946 a_14620_140# a_14950_140# a_14850_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8947 VDD word5.byte3.tinv2.I a_49620_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8948 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8949 word1.byte1.cgate0.inv1.I word1.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8950 VDD buf_sel7.inv0.O buf_sel7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8951 a_151860_10088# a_151650_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X8952 VSS word3.byte3.tinv5.I a_60420_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8953 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8954 VDD word3.byte3.tinv2.I a_49620_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8955 buf_out9.inv1.O buf_out9.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8956 word7.byte1.dff_1.O word7.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8957 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8958 VDD word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8959 VDD a_141060_5492# a_141020_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8960 VDD a_12180_10088# word7.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8961 a_122080_9548# a_122410_9548# a_122310_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X8962 a_17220_3442# word3.byte4.tinv4.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X8963 word4.byte4.tinv7.O buf_out25.inv0.I a_28020_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8964 VDD word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8965 VDD a_4980_10088# a_4940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8966 VSS a_116040_2356# a_116000_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8967 VSS a_7420_7928# a_6420_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8968 a_54780_190# word1.byte3.cgate0.inv1.O a_54220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8969 a_147940_2776# a_146100_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8970 a_18550_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X8971 buf_in25.inv1.O buf_in25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X8972 VDD a_47020_7928# a_46020_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X8973 VDD a_141060_2356# a_141020_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8974 word2.byte4.tinv7.O buf_out25.inv0.I a_28020_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8975 VDD a_40980_6952# word5.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8976 a_65250_9598# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X8977 buf_in7.inv1.O buf_in7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8978 Do19_buf buf_out20.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8979 VSS a_119640_6952# a_119600_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8980 a_159020_5912# a_158230_5632# a_158850_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X8981 VSS a_14620_11064# a_13620_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X8982 a_53220_9714# word7.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X8983 buf_in31.inv1.O buf_in31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8984 VSS buf_in19.inv0.O buf_in19.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8985 VDD word8.byte2.buf_RE1.I word8.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8986 a_104080_140# word1.byte2.dff_7.CLK a_104310_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X8987 VDD a_40980_3816# word3.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X8988 VSS word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8989 VSS word2.byte3.tinv7.I a_67620_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8990 VSS word8.byte1.tinv5.I a_160500_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8991 VDD word1.byte1.tinv7.I a_167700_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X8992 VSS a_119640_3816# a_119600_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X8993 a_115830_4842# a_115210_5632# a_115720_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X8994 VDD buf_in22.inv0.O buf_in22.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8995 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8996 VSS word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X8997 VSS word1.byte3.inv_and.O a_75720_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X8998 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X8999 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.latch0.I0.ENB a_131700_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9000 a_47250_1090# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9001 a_124680_306# buf_out10.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9002 a_140460_2776# word2.byte1.dff_7.CLK a_139900_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9003 VDD buf_we1.inv1.O word8.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9004 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9005 a_108520_9598# a_106680_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9006 a_115110_7978# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9007 a_40770_1706# word2.byte3.cgate0.inv1.O a_40660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9008 a_101430_190# word1.byte2.dff_7.CLK a_101320_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9009 a_115830_1706# a_115210_2496# a_115720_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9010 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9011 word2.byte3.dff_3.O word2.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9012 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9013 VDD a_126840_10088# word7.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9014 word5.gt_re0.OUT buf_sel5.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9015 a_75360_1092# word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9016 a_100810_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9017 VDD a_155460_680# a_155420_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9018 a_56820_9714# word7.byte3.tinv4.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9019 a_11970_7978# word6.byte4.cgate0.inv1.O a_11860_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9020 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.latch0.I0.ENB a_131700_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9021 a_104640_7978# a_104410_8768# a_104080_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9022 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9023 VDD word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9024 word6.byte4.dff_6.O word6.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9025 VSS buf_in15.inv0.I buf_in15.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9026 word5.byte2.dff_6.O word5.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9027 a_20820_3442# word3.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9028 word3.gt_re0.OUT buf_sel3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9029 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9030 word4.byte3.tinv7.O buf_out19.inv0.I a_60420_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9031 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9032 word3.byte2.dff_6.O word3.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9033 VDD word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9034 a_12140_9048# a_11350_8768# a_11970_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9035 word1.byte4.dff_1.O word1.byte4.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9036 a_151860_5492# a_151650_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9037 buf_re.inv1.O buf_re.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9038 a_119040_11114# a_118810_11904# a_118480_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9039 a_58660_4842# a_56820_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9040 buf_in23.inv1.O buf_in23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9041 a_44540_6462# a_43750_6412# a_44370_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9042 word2.byte3.tinv7.O buf_out19.inv0.I a_60420_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9043 Do24_buf buf_out25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9044 a_40940_10498# word7.byte3.cgate0.inv1.O a_40770_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9045 a_25750_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9046 a_155420_7362# word5.byte1.dff_7.CLK a_155250_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9047 a_151540_9048# a_149700_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9048 a_66140_10498# word7.byte3.cgate0.inv1.O a_65970_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9049 VSS a_51780_8628# a_51740_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9050 word1.byte1.dff_5.O word1.byte1.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9051 word2.byte1.tinv7.O word2.byte1.tinv2.EN a_149700_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9052 VSS word2.byte1.buf_RE0.I word2.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9053 a_58660_1706# a_56820_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9054 VDD word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9055 a_44540_3326# a_43750_3276# a_44370_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9056 VDD a_159060_5492# word4.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9057 a_134580_306# word1.byte1.cgate0.nand0.A word1.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9058 a_58980_5492# a_58770_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9059 a_158460_12184# word8.byte1.dff_7.CLK a_157900_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9060 a_155420_4226# word3.byte1.dff_7.CLK a_155250_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9061 a_151030_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9062 VDD buf_out19.inv0.O Do18_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9063 a_118710_11114# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9064 a_162620_11114# word8.byte1.dff_7.CLK a_162450_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9065 a_73020_306# word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9066 a_28020_2660# word2.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9067 VDD a_159060_2356# word2.byte1.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9068 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9069 VDD word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9070 a_58980_2356# a_58770_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9071 VSS buf_sel7.inv0.O buf_sel7.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9072 VDD word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9073 a_126630_190# word1.byte2.dff_7.CLK a_126520_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9074 VDD a_12180_5492# word4.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9075 VSS word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9076 a_144450_11114# a_143830_11904# a_144340_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9077 a_48180_10088# a_47970_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9078 a_90120_9714# word7.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9079 VDD word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9080 a_142500_7976# buf_out8.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9081 a_42420_6578# word5.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9082 VDD a_12180_2356# word2.byte4.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9083 word7.byte4.tinv7.O word7.byte4.tinv4.EN a_17220_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9084 VSS word3.byte1.cgate0.nand0.B a_95160_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9085 a_161830_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9086 a_64020_6578# word5.byte3.tinv6.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9087 word4.byte4.nand.OUT word4.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9088 a_4050_11114# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9089 a_92280_7976# word6.byte2.cgate0.latch0.I0.ENB word6.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9090 a_126800_9598# a_126010_9548# a_126630_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9091 buf_in16.inv1.O buf_in16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9092 VSS a_107680_9548# a_106680_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9093 a_42420_3442# word3.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9094 buf_in9.inv1.O buf_in9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9095 a_117480_11112# word8.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9096 VSS a_44580_10088# word7.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9097 a_150700_11064# word8.byte1.dff_7.CLK a_150930_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9098 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9099 word2.byte4.nand.OUT word2.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9100 buf_in7.inv1.O buf_in7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9101 VDD a_110280_11112# a_111840_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9102 VSS a_144660_11764# a_144620_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9103 buf_in28.inv1.O buf_in28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9104 a_122920_7978# a_121080_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9105 a_65020_6412# a_65350_6412# a_65250_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9106 a_19060_5912# a_17220_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9107 word8.byte1.tinv7.O word8.byte1.tinv0.EN a_142500_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9108 VSS a_46020_1704# a_47580_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9109 buf_in3.inv1.O buf_in3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9110 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9111 a_104410_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9112 a_108800_1090# word1.byte2.dff_7.CLK a_108630_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9113 a_65020_3276# a_65350_3276# a_65250_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9114 VSS buf_in22.inv0.O buf_in22.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9115 VSS a_1380_8628# word6.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9116 VSS a_119640_5492# word4.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9117 VSS a_17220_7976# a_18780_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9118 VDD a_26580_680# word1.byte4.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9119 VSS word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9120 a_158460_5912# word4.byte1.dff_7.CLK a_157900_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9121 a_2820_11112# word8.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9122 VSS a_149700_11112# a_151260_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9123 a_58770_4842# word4.byte3.cgate0.inv1.O a_58660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9124 VSS word8.byte3.tinv4.I a_56820_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9125 a_6420_9714# word7.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9126 a_61750_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9127 a_60420_1704# word2.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9128 a_114880_4792# word4.byte2.dff_7.CLK a_115110_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9129 word8.byte1.tinv7.O buf_out4.inv0.I a_156900_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9130 a_160500_306# word1.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9131 VDD word8.byte4.buf_RE0.O word8.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9132 VSS a_100380_6462# a_101040_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9133 VSS word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9134 VSS word4.byte4.buf_RE0.O word4.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9135 VSS a_144660_680# a_144620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9136 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9137 word8.gt_re1.O word8.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9138 word6.byte1.cgate0.nand0.A word6.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9139 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9140 a_61750_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9141 VDD word4.byte1.tinv6.I a_164100_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9142 VDD buf_sel8.inv0.O buf_sel8.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9143 a_15570_7978# a_14950_8768# a_15460_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9144 a_119640_10088# a_119430_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9145 a_114880_1656# word2.byte2.dff_7.CLK a_115110_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9146 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9147 VSS a_100380_3326# a_101040_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9148 a_134580_6578# word5.byte1.cgate0.nand0.A word5.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9149 word6.byte4.dff_7.O word6.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9150 word7.byte3.tinv7.O word7.byte3.tinv2.EN a_49620_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9151 VDD word2.byte1.tinv6.I a_164100_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9152 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9153 word6.byte2.cgate0.inv1.I word6.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9154 VDD a_153300_7976# a_154860_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9155 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9156 VDD a_166260_5492# a_166220_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9157 a_111610_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9158 word8.byte1.nand.OUT buf_we4.inv1.O a_129540_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9159 a_140850_9598# word7.byte1.dff_7.CLK a_140740_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9160 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9161 buf_in15.inv1.O buf_in15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9162 VDD word6.byte3.tinv3.I a_53220_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9163 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9164 VDD a_166260_2356# a_166220_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9165 a_111610_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9166 Do24_buf buf_out25.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9167 buf_in6.inv1.O buf_in6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9168 a_22770_190# word1.byte4.cgate0.inv1.O a_22660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9169 a_101640_680# a_101430_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9170 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9171 a_4770_4842# a_4150_5632# a_4660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9172 VSS a_151860_11764# word8.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9173 VSS word8.byte2.tinv5.I a_121080_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9174 a_155140_7978# a_153300_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9175 VSS a_8580_680# word1.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9176 VDD a_55380_8628# a_55340_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9177 word6.byte1.buf_RE0.I word6.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9178 VSS word4.byte1.tinv0.I a_142500_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9179 a_26260_2776# a_24420_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9180 a_4770_1706# a_4150_2496# a_4660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9181 VSS word6.byte2.buf_RE1.I word6.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9182 a_55170_6462# a_54550_6412# a_55060_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9183 a_82020_306# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9184 VDD a_122080_140# a_121080_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9185 a_4050_2776# buf_in31.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9186 VSS a_49620_7976# a_51180_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9187 VSS word4.byte2.inv_and.O a_92280_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9188 a_58940_11114# word8.byte3.cgate0.inv1.O a_58770_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9189 word5.byte3.dff_7.O word5.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9190 word6.byte3.tinv7.O word6.byte3.tinv4.EN a_56820_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9191 a_165660_2776# word2.byte1.dff_7.CLK a_165100_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9192 a_55170_3326# a_54550_3276# a_55060_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9193 a_65970_1706# word2.byte3.cgate0.inv1.O a_65860_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9194 word5.byte1.tinv7.O buf_out4.inv0.I a_156900_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9195 VSS buf_sel3.inv0.O buf_sel3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9196 VDD word5.byte2.tinv0.I a_103080_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9197 a_26580_2356# a_26370_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9198 word3.byte3.dff_7.O word3.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9199 a_22050_12184# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9200 word6.byte2.dff_4.O word6.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9201 word3.byte1.tinv7.O buf_out4.inv0.I a_156900_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9202 VDD a_143500_4792# a_142500_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9203 a_25980_4842# a_25750_5632# a_25420_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9204 VSS word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9205 a_47250_12184# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9206 a_4380_190# word1.byte4.cgate0.inv1.O a_3820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9207 VDD word3.byte2.tinv0.I a_103080_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9208 a_160500_11112# buf_out3.inv0.I word8.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9209 a_65580_11114# a_65350_11904# a_65020_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9210 VDD word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9211 a_119040_10498# a_118810_9548# a_118480_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9212 a_46020_3442# word3.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9213 a_161730_6462# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9214 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9215 a_66140_2776# a_65350_2496# a_65970_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9216 VDD a_22980_6952# a_22940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9217 VDD a_143500_1656# a_142500_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9218 a_25980_1706# a_25750_2496# a_25420_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9219 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9220 a_161730_3326# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9221 a_47020_11064# word8.byte3.cgate0.inv1.O a_47250_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9222 VSS a_101640_2356# a_101600_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9223 a_47970_190# word1.byte3.cgate0.inv1.O a_47860_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9224 VDD a_22980_3816# a_22940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9225 a_13620_7976# word6.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9226 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9227 a_65860_12184# a_64020_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9228 a_50850_9598# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9229 Do7_buf buf_out8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9230 a_107910_7362# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9231 a_123200_11114# word8.byte2.dff_7.CLK a_123030_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9232 a_118710_10498# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9233 a_162620_10498# word7.byte1.dff_7.CLK a_162450_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9234 VSS a_119640_680# word1.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9235 VSS word2.byte2.tinv5.I a_121080_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9236 VDD word7.byte4.cgate0.nand0.A word7.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9237 a_107910_4226# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9238 VSS a_46020_11112# a_47580_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9239 VDD buf_in18.inv0.O buf_in18.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9240 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9241 a_144450_9598# a_143830_9548# a_144340_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9242 VDD a_51780_11764# a_51740_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9243 VSS word7.byte1.tinv3.I a_153300_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9244 a_119600_4842# word4.byte2.dff_7.CLK a_119430_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9245 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9246 a_2820_4840# word4.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9247 a_100710_7978# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9248 a_62260_6462# a_60420_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9249 VSS a_122080_1656# a_121080_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9250 a_4380_12184# word8.byte4.cgate0.inv1.O a_3820_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9251 word4.byte3.tinv7.O word4.byte3.tinv6.EN a_64020_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9252 a_122410_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9253 a_110280_9714# word7.byte2.tinv2.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9254 a_4050_10498# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9255 VDD buf_sel4.inv0.O buf_sel4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9256 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9257 a_119600_1706# word2.byte2.dff_7.CLK a_119430_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9258 a_105240_11764# a_105030_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9259 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9260 a_2820_1704# word2.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9261 a_167700_7976# buf_out1.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9262 a_67620_7364# word5.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9263 VDD a_220_140# a_120_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9264 a_62260_3326# a_60420_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9265 a_39820_4792# a_40150_5632# a_40050_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9266 VSS buf_sel5.inv0.I buf_sel5.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9267 VDD word7.byte2.inv_and.O a_92280_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9268 a_150700_9548# word7.byte1.dff_7.CLK a_150930_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9269 a_158230_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9270 buf_in15.inv1.O buf_in15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9271 VSS a_162660_6952# word5.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9272 VSS a_105240_11764# a_105200_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9273 VDD a_110280_9714# a_111840_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9274 a_35760_6578# word5.byte1.cgate0.nand0.B word5.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9275 a_11350_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9276 a_14620_1656# a_14950_2496# a_14850_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9277 VDD word4.byte3.inv_and.O a_75720_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9278 a_24420_6578# buf_out26.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9279 a_62580_6952# a_62370_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9280 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9281 VSS word3.byte3.nand.OUT word3.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9282 a_67620_4228# word3.byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9283 VDD a_139900_6412# a_139800_6462# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9284 a_57820_7928# a_58150_8768# a_58050_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9285 a_75720_7976# word6.byte3.cgate0.latch0.I0.ENB word6.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9286 VSS a_162660_3816# word3.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9287 VDD word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9288 VDD word2.byte3.inv_and.O a_75720_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9289 a_139900_9548# a_140230_9548# a_140130_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9290 a_62580_3816# a_62370_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9291 a_24420_3442# buf_out26.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9292 a_450_7978# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9293 VDD a_139900_3276# a_139800_3326# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9294 buf_in11.inv0.O buf_in11.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9295 buf_in25.inv1.O buf_in25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9296 VDD a_108840_6952# word5.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9297 a_141020_7362# word5.byte1.dff_7.CLK a_140850_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9298 a_117480_7976# word6.byte2.tinv4.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9299 VSS buf_in21.inv0.O buf_in21.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9300 a_46020_9714# word7.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9301 buf_in2.inv0.O Di1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9302 word8.byte2.tinv7.O buf_out12.inv0.I a_117480_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9303 a_155460_8628# a_155250_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9304 word2.byte1.dff_7.CLK word2.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9305 a_54550_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9306 VSS word6.buf_ck1.I word6.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9307 a_141020_4226# word3.byte1.dff_7.CLK a_140850_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9308 VDD a_108840_3816# word3.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9309 VDD buf_in24.inv0.O buf_in24.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9310 a_42420_11112# word8.byte3.tinv0.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9311 VDD buf_in17.inv0.O buf_in17.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9312 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9313 VSS word2.byte1.buf_RE0.I word2.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9314 word4.byte1.cgate0.inv1.I word4.byte1.cgate0.nand0.A a_134580_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9315 word7.byte3.nand.OUT word7.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9316 VSS a_124680_6578# a_126240_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9317 VDD a_101640_8628# word6.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9318 a_42420_1704# word2.byte3.tinv0.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9319 VSS word3.byte2.tinv1.I a_106680_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9320 a_108630_1706# word2.byte2.dff_7.CLK a_108520_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9321 VSS word5.byte1.tinv5.I a_160500_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9322 a_142500_306# buf_out8.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9323 VSS a_26580_10088# a_26540_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9324 VSS a_124680_3442# a_126240_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9325 word8.byte4.tinv7.O buf_out32.inv0.I a_2820_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9326 a_25750_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9327 a_56820_11112# buf_out20.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9328 a_92280_1092# word1.byte2.cgate0.latch0.I0.ENB word1.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9329 a_78780_306# buf_we2.inv1.O word1.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9330 VSS word7.byte3.cgate0.nand0.A a_75360_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9331 a_49620_306# word1.byte3.tinv2.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9332 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9333 word5.byte2.tinv7.O word5.byte2.tinv4.EN a_117480_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9334 VSS a_119640_5492# a_119600_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9335 VSS word5.byte1.nand.OUT word5.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9336 a_166050_9598# word7.byte1.dff_7.CLK a_165940_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9337 buf_out15.inv1.O buf_out15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9338 VSS a_112440_11764# word8.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9339 VSS a_61420_6412# a_60420_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9340 a_36120_4840# word4.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9341 word5.byte1.dff_0.O word5.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9342 VDD buf_in32.inv0.O buf_in32.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9343 word6.byte2.inv_and.O word6.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9344 VDD a_20820_6578# a_22380_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9345 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9346 a_110280_9714# word7.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9347 a_126840_680# a_126630_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9348 Do5_buf buf_out6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9349 word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.latch0.I0.ENB a_36120_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9350 a_50620_6412# a_50950_6412# a_50850_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9351 a_36120_1704# word2.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9352 word3.byte1.dff_0.O word3.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9353 VSS a_61420_3276# a_60420_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9354 buf_re.inv1.O buf_re.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9355 VDD a_20820_3442# a_22380_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9356 VSS word8.byte4.buf_RE0.O word8.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9357 a_161500_6412# word5.byte1.dff_7.CLK a_161730_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9358 a_58940_10498# word7.byte3.cgate0.inv1.O a_58770_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9359 VSS word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9360 VSS word4.byte1.tinv7.I a_167700_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9361 a_148050_190# a_147430_140# a_147940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9362 a_50620_3276# a_50950_3276# a_50850_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9363 VDD a_13620_11112# a_15180_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9364 VSS word6.gt_re0.OUT word6.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9365 a_161500_3276# word3.byte1.dff_7.CLK a_161730_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9366 a_124680_4840# word4.byte2.tinv6.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9367 VDD a_104080_11064# a_103080_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9368 VDD buf_in1.inv0.O buf_in1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9369 VSS a_4980_11764# word8.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9370 word4.byte2.dff_6.O word4.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9371 a_33420_2660# word2.byte4.cgate0.nand0.A word2.byte4.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9372 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9373 a_75360_5796# word4.byte1.cgate0.nand0.B word4.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9374 VDD word5.byte2.tinv7.I a_128280_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9375 a_100480_4792# word4.byte2.dff_7.CLK a_100710_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9376 a_65580_10498# a_65350_9548# a_65020_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9377 word1.byte1.cgate0.nand0.A word1.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9378 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9379 VSS word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9380 dec8.and4_4.nand1.OUT A2 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9381 word8.buf_sel0.O buf_sel8.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9382 word1.byte4.dff_3.O word1.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9383 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9384 a_154530_9048# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9385 a_100480_1656# word2.byte2.dff_7.CLK a_100710_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9386 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9387 VDD word3.byte2.tinv7.I a_128280_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9388 a_143730_12184# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9389 a_149700_4840# word4.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9390 a_44540_5912# a_43750_5632# a_44370_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9391 a_15570_11114# word8.byte4.cgate0.inv1.O a_15460_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9392 VSS a_40980_680# word1.byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9393 word1.byte2.cgate0.inv1.I word1.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9394 a_43650_4842# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9395 a_35760_11112# word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9396 a_47020_9548# word7.byte3.cgate0.inv1.O a_47250_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9397 VDD a_116040_6952# a_116000_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9398 VDD a_139800_190# a_140460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9399 a_112230_7978# word6.byte2.dff_7.CLK a_112120_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9400 word4.byte2.tinv7.O buf_out15.inv0.I a_106680_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9401 a_147940_7362# a_146100_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9402 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9403 VDD word4.byte2.buf_RE1.I word4.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9404 word6.byte1.tinv7.O buf_out3.inv0.I a_160500_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9405 VDD word1.byte3.tinv3.I a_53220_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9406 VDD a_151860_5492# a_151820_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9407 a_149700_1704# word2.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9408 a_28020_3442# word3.byte4.tinv7.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9409 buf_in11.inv1.O buf_in11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9410 a_43650_1706# buf_in23.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9411 word5.gt_re1.O word5.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9412 VDD a_116040_3816# a_116000_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9413 a_143500_11064# word8.byte1.dff_7.CLK a_143730_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9414 VSS a_126840_2356# a_126800_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9415 a_123200_10498# word7.byte2.dff_7.CLK a_123030_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9416 a_104920_190# a_103080_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9417 a_147940_4226# a_146100_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9418 a_144620_9598# a_143830_9548# a_144450_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9419 word2.byte2.tinv7.O buf_out15.inv0.I a_106680_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9420 VDD word2.byte2.buf_RE1.I word2.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9421 VDD a_57820_7928# a_56820_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9422 VSS word5.byte4.tinv7.I a_28020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9423 VDD a_151860_2356# a_151820_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9424 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9425 VDD a_21820_9548# a_20820_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9426 a_220_4792# word4.byte4.cgate0.inv1.O a_450_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9427 VSS word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9428 VDD buf_out14.inv0.O buf_out14.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9429 VDD a_47020_9548# a_46020_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9430 VDD Di27 buf_in28.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9431 a_140740_7978# a_139800_7978# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9432 VDD a_51780_10088# a_51740_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9433 VDD a_40980_8628# a_40940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9434 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9435 a_153300_7976# word6.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9436 a_6420_9714# buf_out31.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9437 a_159060_8628# a_158850_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9438 VSS buf_in17.inv0.O buf_in17.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9439 VSS buf_out5.inv0.O Do4_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9440 a_140460_7362# a_140230_6412# a_139900_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9441 a_11860_2776# a_10020_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9442 a_220_1656# word2.byte4.cgate0.inv1.O a_450_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9443 a_58150_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9444 a_40770_6462# a_40150_6412# a_40660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9445 a_780_11114# a_550_11904# a_220_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9446 word8.byte4.cgate0.inv1.I word8.byte4.cgate0.nand0.A a_33420_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9447 word5.byte3.dff_3.O word5.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9448 a_55060_9048# a_53220_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9449 a_105240_10088# a_105030_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9450 a_140460_4226# a_140230_3276# a_139900_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9451 a_40770_3326# a_40150_3276# a_40660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9452 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9453 a_125910_7978# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9454 a_58050_1090# buf_in19.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9455 buf_in19.inv1.O buf_in19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9456 VSS word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9457 a_115440_1090# a_115210_140# a_114880_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9458 a_12180_2356# a_11970_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9459 word3.byte3.dff_3.O word3.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9460 word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.latch0.I0.ENB a_92280_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9461 a_155460_680# a_155250_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9462 word6.byte2.dff_0.O word6.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9463 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9464 VSS a_155460_8628# word6.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9465 a_65020_4792# a_65350_5632# a_65250_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9466 a_107680_1656# a_108010_2496# a_107910_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9467 word3.byte2.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9468 buf_sel6.inv1.O buf_sel6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9469 word5.byte4.inv_and.O word5.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9470 VSS a_24420_9714# a_25980_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9471 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9472 word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.latch0.I0.ENB a_92280_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9473 a_51740_2776# a_50950_2496# a_51570_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9474 a_92280_12068# word8.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9475 a_60420_3442# word3.byte3.tinv5.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9476 word3.byte4.inv_and.O word3.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9477 a_25750_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9478 VSS word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9479 a_13620_306# word1.byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9480 VDD word4.byte3.cgate0.inv1.I word4.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9481 word8.byte3.cgate0.inv1.I word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9482 a_21820_7928# word6.byte4.cgate0.inv1.O a_22050_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9483 a_165100_9548# a_165430_9548# a_165330_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9484 a_22940_9048# a_22150_8768# a_22770_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9485 a_123200_6462# a_122410_6412# a_123030_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9486 a_125680_140# a_126010_140# a_125910_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9487 VSS a_104080_6412# a_103080_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9488 buf_in8.inv1.O buf_in8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9489 a_61750_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9490 VDD word4.byte4.tinv4.I a_17220_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9491 VSS a_159060_2356# a_159020_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9492 a_104410_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9493 VDD word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9494 VDD word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9495 VDD buf_in10.inv0.O buf_in10.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9496 a_25750_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9497 VSS word8.byte1.buf_RE1.I word8.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9498 a_123200_3326# a_122410_3276# a_123030_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9499 VSS a_100380_4842# a_101040_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9500 a_4940_1090# word1.byte4.cgate0.inv1.O a_4770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9501 VSS a_104080_3276# a_103080_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9502 a_61980_190# word1.byte3.cgate0.inv1.O a_61420_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9503 VDD word2.byte4.tinv4.I a_17220_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9504 a_167700_10500# word7.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9505 VSS buf_in1.inv0.O buf_in1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9506 VDD word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9507 VDD a_19380_5492# a_19340_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9508 VSS buf_in23.inv0.O buf_in23.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9509 a_106680_1704# word2.byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9510 VSS word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9511 a_161830_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9512 a_147100_140# word1.byte1.dff_7.CLK a_147330_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9513 a_160500_4840# word4.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9514 buf_in30.inv1.O buf_in30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9515 VSS a_117480_7976# a_119040_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9516 word2.byte4.dff_2.O word2.byte4.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9517 VDD a_19380_2356# a_19340_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9518 a_158850_4842# a_158230_5632# a_158740_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9519 dec8.and4_6.nand0.A A0 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9520 a_25750_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9521 VDD a_126840_8628# word6.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9522 VDD a_22980_5492# word4.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9523 VSS word7.byte1.buf_RE1.I word7.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9524 a_67620_2660# word2.byte3.tinv7.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9525 a_167700_1092# buf_out1.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9526 a_78780_12068# buf_we2.inv1.O word8.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9527 VDD buf_sel3.inv0.O buf_sel3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9528 a_158130_7978# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9529 a_121080_6578# word5.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9530 a_158850_1706# a_158230_2496# a_158740_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9531 VSS word1.gt_re1.O word1.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9532 a_40050_12184# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9533 VDD a_22980_2356# word2.byte4.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9534 word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.latch0.I0.O a_132960_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9535 a_143830_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9536 word4.byte1.inv_and.O word4.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9537 a_147430_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9538 a_121080_3442# word3.byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9539 a_10020_6578# buf_out30.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9540 a_75720_1092# word1.byte3.cgate0.latch0.I0.ENB word1.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9541 word5.byte1.dff_7.O word5.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9542 word2.byte1.inv_and.O word2.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9543 a_18780_2776# word2.byte4.cgate0.inv1.O a_18220_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9544 word3.byte1.cgate0.latch0.I0.O word3.byte1.cgate0.latch0.I0.O a_132960_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9545 VDD a_46020_6578# a_47580_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9546 VDD a_149700_4840# a_151260_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9547 a_43420_7928# a_43750_8768# a_43650_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9548 a_11250_2776# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9549 VSS buf_out14.inv0.I buf_out14.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9550 VSS a_142500_306# a_144060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9551 VSS a_8580_8628# a_8540_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9552 word3.byte4.tinv7.O word3.byte4.tinv5.EN a_20820_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9553 a_10020_3442# buf_out30.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9554 word6.byte3.cgate0.inv1.I word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9555 word3.byte1.dff_7.O word3.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9556 a_50850_11114# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9557 a_104640_12184# word8.byte2.dff_7.CLK a_104080_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9558 VDD a_13620_9714# a_15180_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9559 a_144060_9598# word7.byte1.dff_7.CLK a_143500_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9560 VDD a_149700_1704# a_151260_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9561 VDD a_46020_3442# a_47580_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9562 a_116000_11114# word8.byte2.dff_7.CLK a_115830_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9563 a_44370_9598# word7.byte3.cgate0.inv1.O a_44260_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9564 word6.byte4.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9565 a_103080_7976# word6.byte2.tinv0.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9566 a_14850_6462# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9567 word7.byte3.dff_4.O word7.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9568 VSS buf_in7.inv0.O buf_in7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9569 VSS buf_out20.inv0.O Do19_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9570 VDD a_39720_7978# a_40380_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9571 VDD a_39820_11064# a_39720_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9572 VDD buf_out1.inv0.O Do0_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9573 a_14850_3326# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9574 a_161730_5912# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9575 a_104310_12184# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9576 VDD word7.byte1.cgate0.nand0.B word7.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9577 dec8.and4_6.nand1.OUT A2 a_75360_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9578 a_1170_7978# word6.byte4.cgate0.inv1.O a_1060_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9579 VSS a_110280_6578# a_111840_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9580 a_26370_190# a_25750_140# a_26260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9581 a_142500_306# word1.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9582 VSS word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9583 word6.byte2.dff_1.O word6.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9584 word2.byte4.tinv7.O word2.byte4.tinv7.EN a_28020_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9585 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9586 a_104080_11064# word8.byte2.dff_7.CLK a_104310_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9587 a_143500_9548# word7.byte1.dff_7.CLK a_143730_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9588 VSS a_110280_3442# a_111840_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9589 VDD word5.byte3.cgate0.nand0.A word5.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9590 VDD a_164100_306# a_165660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9591 a_126240_4842# a_126010_5632# a_125680_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9592 VSS a_47020_4792# a_46020_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9593 a_95160_6578# word5.byte2.cgate0.nand0.A word5.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9594 word5.byte2.tinv7.O word5.byte2.tinv0.EN a_103080_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9595 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9596 word1.byte2.inv_and.O word1.byte2.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9597 buf_sel5.inv1.O buf_sel5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9598 word8.byte1.dff_4.O word8.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9599 word5.byte4.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9600 buf_in15.inv1.O buf_in15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9601 VDD word3.byte3.cgate0.nand0.A word3.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9602 a_51180_2776# word2.byte3.cgate0.inv1.O a_50620_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9603 VDD word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9604 a_64020_11112# word8.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9605 a_26540_7978# word6.byte4.cgate0.inv1.O a_26370_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9606 word5.byte3.tinv7.O buf_out24.inv0.I a_42420_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9607 word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.latch0.I0.ENB a_36120_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9608 a_126240_1706# a_126010_2496# a_125680_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9609 VDD word8.buf_sel0.O word8.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9610 a_112440_680# a_112230_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9611 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9612 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9613 VSS buf_out13.inv0.O buf_out13.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9614 a_26260_7362# a_24420_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9615 a_780_10498# a_550_9548# a_220_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9616 a_22380_9048# word6.byte4.cgate0.inv1.O a_21820_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9617 a_4050_7362# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9618 VDD a_66180_680# a_66140_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9619 VDD a_143500_9548# a_142500_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9620 VDD word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9621 buf_in27.inv1.O buf_in27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9622 buf_in13.inv0.O buf_in13.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9623 word3.byte3.tinv7.O buf_out24.inv0.I a_42420_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9624 a_165940_7978# a_164100_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9625 a_62260_5912# a_60420_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9626 a_54780_6462# word5.byte3.cgate0.inv1.O a_54220_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9627 VDD word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9628 VSS word1.byte3.buf_RE0.O word1.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9629 buf_in4.inv0.O Di3 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9630 a_26260_4226# a_24420_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9631 VSS buf_out27.inv0.O Do26_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9632 VSS a_8580_11764# a_8540_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9633 a_4050_4226# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9634 a_165660_7362# a_165430_6412# a_165100_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9635 a_65970_6462# a_65350_6412# a_65860_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9636 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9637 a_4380_1090# a_4150_140# a_3820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9638 a_26580_6952# a_26370_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9639 a_54780_3326# word3.byte3.cgate0.inv1.O a_54220_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9640 VDD buf_out30.inv0.I buf_out30.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X9641 word8.byte4.tinv7.O word8.byte4.tinv1.EN a_6420_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9642 VSS a_162660_5492# word4.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9643 a_165660_4226# a_165430_3276# a_165100_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9644 a_62580_5492# a_62370_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9645 a_111610_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9646 a_65970_3326# a_65350_3276# a_65860_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9647 VDD word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9648 Do18_buf buf_out19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9649 a_167700_306# word1.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9650 a_26580_3816# a_26370_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9651 word7.byte4.tinv7.O word7.byte4.tinv1.EN a_6420_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9652 a_157900_4792# word4.byte1.dff_7.CLK a_158130_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9653 a_77700_13636# dec8.and4_7.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9654 a_66140_7362# word5.byte3.cgate0.inv1.O a_65970_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9655 word6.byte2.dff_7.O word6.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9656 word2.byte3.tinv7.O word2.byte3.tinv5.EN a_60420_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9657 a_124680_3442# word3.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9658 a_108840_6952# a_108630_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9659 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9660 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9661 word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.latch0.I0.ENB a_75720_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9662 VDD word8.byte1.cgate0.nand0.B word8.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9663 a_162660_10088# a_162450_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9664 VDD a_101640_6952# a_101600_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9665 word1.byte1.tinv7.O buf_out3.inv0.I a_160500_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9666 a_157900_1656# word2.byte1.dff_7.CLK a_158130_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9667 VSS a_151860_680# a_151820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9668 VSS word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9669 VSS word7.byte3.buf_RE0.O word7.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9670 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9671 word3.byte3.cgate0.nand0.A word3.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9672 a_66140_4226# word3.byte3.cgate0.inv1.O a_65970_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9673 word6.byte1.cgate0.inv1.I word6.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9674 word5.byte4.cgate0.inv1.I word5.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9675 a_108840_3816# a_108630_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9676 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9677 word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.latch0.I0.ENB a_75720_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9678 VDD a_101640_3816# a_101600_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9679 word3.byte4.cgate0.inv1.O word3.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9680 a_47020_7928# word6.byte3.cgate0.inv1.O a_47250_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9681 a_154630_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9682 VDD word6.gt_re1.O word6.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9683 VSS word1.byte2.tinv3.I a_113880_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9684 a_128280_10500# word7.byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9685 VSS word5.byte4.tinv3.I a_13620_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9686 VSS a_66180_6952# word5.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9687 word3.byte4.cgate0.inv1.I word3.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9688 VSS buf_in9.inv0.O buf_in9.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9689 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9690 VSS a_6420_7976# a_7980_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9691 a_144660_680# a_144450_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9692 a_154630_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9693 VSS a_124680_4840# a_126240_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9694 a_53220_7976# buf_out21.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9695 VSS a_66180_3816# word3.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9696 a_43750_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9697 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9698 Do29_buf buf_out30.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9699 VDD buf_in26.inv0.O buf_in26.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9700 VSS word8.byte1.nand.B a_39180_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9701 a_111510_1090# buf_in13.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9702 a_40660_9048# a_39720_7978# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9703 word6.buf_sel0.O buf_sel6.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9704 VDD a_25420_6412# a_24420_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9705 a_44540_12184# a_43750_11904# a_44370_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9706 a_113880_11112# buf_out13.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9707 VDD word7.byte3.tinv7.I a_67620_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9708 VSS word3.byte4.dff_0.O_bar a_2820_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9709 a_142500_4840# word4.byte1.tinv0.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9710 a_65820_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9711 word4.byte1.dff_0.O word4.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9712 a_108010_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9713 a_147430_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9714 a_121080_9714# word7.byte2.tinv5.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9715 VSS word6.byte3.tinv1.I a_46020_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9716 a_57820_140# a_58150_140# a_58050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9717 VSS word2.byte1.nand.B a_39180_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9718 a_14620_6412# word5.byte4.cgate0.inv1.O a_14850_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9719 a_101040_1090# a_100810_140# a_100480_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9720 VDD buf_in32.inv0.O buf_in32.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9721 VDD buf_sel4.inv0.O buf_sel4.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9722 VDD a_25420_3276# a_24420_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9723 a_92280_5796# word4.byte2.cgate0.latch0.I0.O word4.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9724 VDD word5.byte1.tinv1.I a_146100_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9725 VSS word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9726 VSS a_141060_8628# word6.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9727 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9728 a_50620_4792# a_50950_5632# a_50850_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9729 a_93540_10500# word7.byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9730 a_40980_8628# a_40770_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9731 a_14620_3276# word3.byte4.cgate0.inv1.O a_14850_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9732 VSS a_10020_9714# a_11580_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9733 word7.gt_re3.I word7.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9734 VDD word3.byte1.tinv1.I a_146100_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9735 a_51180_12184# word8.byte3.cgate0.inv1.O a_50620_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9736 VSS a_161500_9548# a_160500_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9737 word4.byte3.dff_2.O word4.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9738 a_50850_10498# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9739 word3.byte1.nand.B word3.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9740 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9741 a_7650_9598# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9742 a_116000_10498# word7.byte2.dff_7.CLK a_115830_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9743 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9744 VDD word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9745 word8.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9746 VSS word1.byte1.buf_RE1.I word1.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9747 word3.byte3.tinv7.O word3.byte3.tinv1.EN a_46020_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9748 a_162450_6462# word5.byte1.dff_7.CLK a_162340_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9749 word2.byte3.dff_2.O word2.byte3.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9750 VSS a_144660_2356# a_144620_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9751 a_44370_11114# a_43750_11904# a_44260_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9752 VDD a_39820_9548# a_39720_9598# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9753 VDD buf_out9.inv0.O buf_out9.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9754 a_162450_3326# word3.byte1.dff_7.CLK a_162340_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9755 a_40050_6462# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9756 VDD a_143500_140# a_142500_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9757 a_123240_5492# a_123030_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9758 buf_we4.inv1.O buf_we4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9759 VSS buf_out24.inv0.I buf_out24.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9760 word6.byte4.tinv7.O buf_out29.inv0.I a_13620_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9761 VDD a_64020_7976# a_65580_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9762 a_1060_11114# a_120_11114# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9763 VSS word6.byte1.nand.B a_78780_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9764 VSS word2.byte1.tinv6.I a_164100_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9765 word4.byte1.cgate0.nand0.A word4.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9766 a_40050_3326# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9767 VSS word8.byte4.tinv2.I a_10020_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9768 a_62580_11764# a_62370_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9769 a_108630_6462# a_108010_6412# a_108520_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9770 VSS a_103080_7976# a_104640_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9771 VDD a_112440_680# word1.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9772 a_123240_2356# a_123030_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9773 buf_in21.inv1.O buf_in21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9774 a_104080_9548# word7.byte2.dff_7.CLK a_104310_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9775 a_108630_3326# a_108010_3276# a_108520_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9776 word4.byte2.cgate0.inv1.I word4.byte2.cgate0.nand0.A a_95160_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9777 VSS a_105240_10088# a_105200_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9778 word8.byte3.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9779 word8.byte2.dff_4.O word8.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9780 word7.byte1.dff_4.O word7.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9781 VSS a_25420_7928# a_24420_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9782 a_143730_7978# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9783 a_153300_9714# word7.byte1.tinv3.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9784 VSS word4.byte3.tinv3.I a_53220_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9785 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9786 VDD word8.byte4.tinv6.I a_24420_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9787 a_101430_7978# a_100810_8768# a_101320_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9788 word4.byte4.tinv7.O buf_out32.inv0.I a_2820_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9789 word5.byte2.tinv7.O word5.byte2.tinv7.EN a_128280_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9790 buf_sel6.inv1.O buf_sel6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9791 word5.byte1.dff_3.O word5.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9792 word3.byte2.buf_RE1.I word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9793 word5.byte3.tinv7.O buf_out17.inv0.I a_67620_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9794 a_78780_6578# buf_we2.inv1.O word5.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9795 VSS word5.byte2.nand.OUT word5.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9796 word2.byte4.tinv7.O buf_out32.inv0.I a_2820_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9797 word1.byte3.cgate0.inv1.I word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9798 word8.byte3.tinv7.O buf_out22.inv0.I a_49620_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9799 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9800 buf_in12.inv0.O buf_in12.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9801 a_36120_6578# word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9802 VDD word4.byte1.cgate0.nand0.B word4.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9803 word3.byte1.dff_3.O word3.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9804 a_47580_9048# word6.byte3.cgate0.inv1.O a_47020_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9805 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9806 word8.byte4.dff_0.O word8.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9807 VSS word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9808 word3.byte3.tinv7.O buf_out17.inv0.I a_67620_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9809 VDD a_54220_4792# a_53220_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9810 buf_in32.inv1.O buf_in32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9811 VDD word2.byte1.cgate0.nand0.B word2.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9812 word7.byte3.dff_0.O word7.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9813 VSS buf_out8.inv0.O Do7_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9814 VSS buf_out29.inv0.I buf_out29.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9815 VDD a_54220_1656# a_53220_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9816 VDD buf_in1.inv0.O buf_in1.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9817 a_156900_11112# word8.byte1.tinv4.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9818 a_112120_2776# a_110280_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9819 buf_in23.inv0.O Di22 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9820 a_12140_11114# word8.byte4.cgate0.inv1.O a_11970_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9821 a_44260_7978# a_42420_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9822 a_18220_9548# a_18550_9548# a_18450_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9823 VSS a_143500_1656# a_142500_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9824 buf_in32.inv0.O Di31 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9825 a_11970_190# a_11350_140# a_11860_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9826 VSS word6.buf_ck1.I word6.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9827 word1.byte4.dff_6.O word1.byte4.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9828 a_123200_5912# a_122410_5632# a_123030_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9829 VSS a_51780_11764# word8.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9830 VDD a_144660_8628# word6.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9831 a_115720_6462# a_113880_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9832 a_122310_4842# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9833 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9834 a_3820_1656# a_4150_2496# a_4050_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9835 VSS word3.byte1.tinv2.I a_149700_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9836 VSS buf_sel1.inv0.I buf_sel1.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9837 word7.gt_re3.I word7.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9838 a_44580_8628# a_44370_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9839 VDD a_126840_6952# a_126800_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9840 VSS a_15780_2356# word2.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9841 a_123030_7978# word6.byte2.dff_7.CLK a_122920_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9842 a_14950_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9843 a_106680_3442# word3.byte2.tinv1.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9844 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9845 a_111840_4842# a_111610_5632# a_111280_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9846 a_13620_4840# word4.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9847 a_11350_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9848 a_122310_1706# buf_in10.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9849 a_115720_3326# a_113880_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9850 VDD dec8.and4_5.nand1.B dec8.and4_4.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9851 word5.byte3.buf_RE0.O word5.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9852 a_12140_1090# word1.byte4.cgate0.inv1.O a_11970_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9853 a_160500_6578# word5.byte1.tinv5.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X9854 VSS word8.buf_ck1.I word8.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9855 a_7420_6412# a_7750_6412# a_7650_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9856 VSS word7.byte3.tinv6.I a_64020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9857 VDD a_126840_3816# a_126800_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9858 a_117480_7976# word6.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9859 word1.byte1.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B a_132960_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9860 a_111840_1706# a_111610_2496# a_111280_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9861 VDD word8.byte3.buf_RE0.O word8.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9862 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9863 VSS word3.byte3.buf_RE0.O word3.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9864 VSS buf_out9.inv0.I buf_out9.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X9865 a_43750_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9866 a_550_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9867 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9868 a_140740_11114# a_139800_11114# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9869 VDD word6.byte1.nand.B word6.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9870 a_151540_1090# a_149700_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9871 VDD a_43420_11064# a_42420_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X9872 a_11860_7362# a_10020_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9873 VSS word1.byte2.buf_RE1.I word1.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9874 a_7420_3276# a_7750_3276# a_7650_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9875 VDD a_51780_680# a_51740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9876 VDD buf_in13.inv0.O buf_in13.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9877 word4.byte4.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9878 VSS a_142500_1704# a_144060_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9879 a_2820_1704# word2.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9880 a_11860_4226# a_10020_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9881 VSS buf_in25.inv0.O buf_in25.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9882 VSS buf_in11.inv0.I buf_in11.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9883 a_108010_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9884 word6.byte2.tinv7.O word6.byte2.tinv5.EN a_121080_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9885 word2.byte4.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9886 a_12180_6952# a_11970_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9887 VDD buf_in7.inv0.O buf_in7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9888 VDD a_106680_7976# a_108240_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9889 a_65860_9048# a_64020_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9890 VSS a_146100_6578# a_147660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9891 a_141020_12184# a_140230_11904# a_140850_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9892 a_167700_5796# word4.byte1.tinv7.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9893 a_166220_12184# a_165430_11904# a_166050_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9894 a_53220_9714# buf_out21.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9895 a_107680_6412# word5.byte2.dff_7.CLK a_107910_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9896 word4.byte1.dff_7.O word4.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9897 VSS buf_in31.inv0.O buf_in31.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9898 buf_in19.inv1.O buf_in19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9899 a_12180_3816# a_11970_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9900 VSS word6.gt_re1.O word6.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9901 VSS word2.byte3.inv_and.O a_75720_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9902 VSS word1.byte3.tinv1.I a_46020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9903 VSS a_146100_3442# a_147660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9904 a_143500_4792# word4.byte1.dff_7.CLK a_143730_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9905 a_67620_12068# word8.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9906 a_51740_7362# word5.byte3.cgate0.inv1.O a_51570_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9907 VDD a_123240_5492# word4.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9908 VDD Di21 buf_in22.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9909 VSS word7.byte2.cgate0.inv1.I word7.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9910 a_107680_3276# word3.byte2.dff_7.CLK a_107910_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9911 a_118480_1656# a_118810_2496# a_118710_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9912 a_75720_5796# word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9913 a_66180_8628# a_65970_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9914 a_128280_7364# buf_out9.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9915 word1.byte1.cgate0.inv1.I word1.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9916 buf_sel2.inv1.O buf_sel2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9917 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9918 VSS a_48180_6952# a_48140_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9919 a_143500_1656# word2.byte1.dff_7.CLK a_143730_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9920 VDD a_123240_2356# word2.byte2.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9921 a_51740_4226# word3.byte3.cgate0.inv1.O a_51570_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9922 a_14850_5912# buf_in28.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9923 a_149700_4840# buf_out6.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9924 VDD buf_sel2.inv0.I buf_sel2.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9925 a_104410_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9926 VDD word1.gt_re1.O word1.gt_re3.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9927 VDD a_159060_6952# a_159020_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9928 a_101600_9048# a_100810_8768# a_101430_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9929 a_155250_7978# word6.byte1.dff_7.CLK a_155140_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9930 a_44370_9598# a_43750_9548# a_44260_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9931 a_128280_4228# buf_out9.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9932 a_7650_12184# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X9933 word8.byte4.dff_5.O word8.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9934 VSS a_19380_8628# word6.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9935 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9936 VSS a_48180_3816# a_48140_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9937 a_148260_11764# a_148050_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X9938 VSS a_114880_6412# a_113880_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9939 VSS word1.gt_re0.OUT word1.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9940 a_24420_9714# word7.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9941 a_149700_1704# buf_out6.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9942 VSS buf_out15.inv0.O buf_out15.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9943 VSS a_51780_6952# word5.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9944 VDD a_159060_3816# a_159020_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9945 a_104410_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9946 VDD word6.byte3.buf_RE0.O word6.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9947 VDD buf_re.inv1.O word6.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9948 buf_in32.inv1.O buf_in32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9949 a_53220_306# buf_out21.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X9950 VSS a_113880_11112# a_115440_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9951 a_1060_10498# a_120_9598# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9952 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X9953 VSS a_110280_4840# a_111840_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X9954 VDD a_1380_680# word1.byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9955 VDD a_17220_306# a_18780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9956 a_7420_11064# word8.byte4.cgate0.inv1.O a_7650_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X9957 VDD a_126840_11764# a_126800_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9958 a_62580_10088# a_62370_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X9959 VSS a_114880_3276# a_113880_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X9960 word5.byte4.dff_2.O word5.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9961 VSS a_51780_3816# word3.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X9962 word7.byte1.cgate0.inv1.I word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9963 VSS buf_re.inv0.O buf_re.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9964 VDD buf_out4.inv0.O Do3_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9965 word3.byte4.dff_2.O word3.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9966 VDD buf_out25.inv0.I buf_out25.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X9967 a_147660_190# word1.byte1.dff_7.CLK a_147100_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9968 word7.byte2.dff_4.O word7.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9969 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9970 VDD a_19380_11764# word8.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X9971 word1.byte3.tinv7.O word1.byte3.tinv0.EN a_42420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9972 word6.byte4.dff_0.O word6.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9973 VDD word5.byte1.inv_and.O a_131700_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9974 a_36120_2660# word2.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9975 a_8540_2776# a_7750_2496# a_8370_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9976 a_18780_7362# a_18550_6412# a_18220_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9977 word4.byte2.inv_and.O word4.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9978 buf_sel8.inv1.O buf_sel8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9979 VDD word8.byte1.tinv1.I a_146100_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9980 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9981 a_126630_7978# a_126010_8768# a_126520_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9982 a_11250_7362# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9983 a_22770_4842# a_22150_5632# a_22660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9984 word6.byte1.dff_1.O word6.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X9985 a_142500_3442# word3.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9986 VDD word3.byte1.inv_and.O a_131700_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9987 a_54780_5912# word4.byte3.cgate0.inv1.O a_54220_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9988 word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.latch0.I0.O a_36120_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9989 word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.latch0.I0.O a_93540_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X9990 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X9991 word7.byte4.dff_0.O word7.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X9992 a_122080_7928# a_122410_8768# a_122310_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X9993 a_18780_4226# a_18550_3276# a_18220_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X9994 a_15460_9598# a_13620_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X9995 a_22770_1706# a_22150_2496# a_22660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X9996 VSS word3.byte2.buf_RE1.I word3.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X9997 a_92280_3442# word3.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X9998 a_11250_4226# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X9999 VDD buf_we1.inv1.O word5.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10000 a_4770_190# word1.byte4.cgate0.inv1.O a_4660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10001 a_22050_2776# buf_in26.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10002 word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.latch0.I0.O a_93540_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10003 VSS word5.byte1.cgate0.nand0.B a_73020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10004 VDD word4.byte3.tinv5.I a_60420_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10005 a_11580_7978# a_11350_8768# a_11020_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10006 a_154860_9598# word7.byte1.dff_7.CLK a_154300_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10007 a_166220_6462# a_165430_6412# a_166050_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10008 VDD buf_in16.inv0.O buf_in16.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10009 a_65250_9048# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10010 a_1060_2776# a_120_1706# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10011 VDD buf_we1.inv1.O word3.byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10012 a_117480_11112# word8.byte2.tinv4.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10013 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10014 VSS word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10015 word1.byte4.tinv7.O buf_out29.inv0.I a_13620_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10016 a_147430_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10017 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10018 a_12140_10498# word7.byte4.cgate0.inv1.O a_11970_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10019 a_15780_10088# a_15570_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10020 VDD a_49620_306# a_51180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10021 word7.byte1.tinv7.O buf_out7.inv0.I a_146100_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10022 VDD word2.byte3.tinv5.I a_60420_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10023 VSS buf_in7.inv0.O buf_in7.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10024 a_17220_4840# buf_out28.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10025 a_166220_3326# a_165430_3276# a_166050_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10026 a_162340_4842# a_160500_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10027 VDD a_62580_5492# a_62540_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10028 a_108840_5492# a_108630_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10029 a_4660_6462# a_2820_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10030 a_149700_1704# word2.byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10031 a_17220_1704# buf_out28.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10032 a_55340_9598# a_54550_9548# a_55170_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10033 a_162340_1706# a_160500_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10034 VDD a_62580_2356# a_62540_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10035 Do21_buf buf_out22.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10036 a_108520_9048# a_106680_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10037 a_10020_6578# word5.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10038 word1.byte2.dff_4.O word1.byte2.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10039 a_4660_3326# a_2820_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10040 word1.byte3.tinv7.O word1.byte3.tinv7.EN a_67620_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10041 word2.byte2.tinv7.O word2.byte2.tinv1.EN a_106680_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10042 VSS word2.byte2.buf_RE1.I word2.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10043 Do2_buf buf_out3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10044 a_2820_11112# word8.byte4.tinv0.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10045 word4.byte1.tinv7.O word4.byte1.tinv5.EN a_160500_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10046 dec8.and4_1.nand1.OUT dec8.and4_3.nand1.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10047 VSS a_66180_5492# word4.byte3.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10048 a_4980_6952# a_4770_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10049 a_108010_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10050 a_132960_3442# word3.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10051 a_10020_3442# word3.byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10052 a_51180_7362# a_50950_6412# a_50620_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10053 a_164100_6578# word5.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10054 a_75360_12850# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10055 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10056 VSS a_57820_4792# a_56820_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10057 a_43980_12184# word8.byte3.cgate0.inv1.O a_43420_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10058 VSS word7.byte1.buf_RE1.I word7.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10059 a_101320_11114# a_100380_11114# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10060 a_140740_10498# a_139800_9598# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10061 a_4980_3816# a_4770_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10062 VSS word8.gt_re1.O word8.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10063 a_105200_7978# word6.byte2.dff_7.CLK a_105030_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10064 buf_we3.inv1.O buf_we3.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10065 word7.byte1.nand.B word7.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10066 a_164100_3442# word3.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10067 a_51180_4226# a_50950_3276# a_50620_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10068 word5.byte3.tinv7.O buf_out21.inv0.I a_53220_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10069 a_61980_2776# word2.byte3.cgate0.inv1.O a_61420_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10070 VDD word8.byte1.buf_RE0.I word8.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10071 a_25420_11064# a_25750_11904# a_25650_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10072 VSS buf_in12.inv0.O buf_in12.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10073 VDD a_165100_11064# a_164100_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10074 word3.byte3.tinv7.O buf_out21.inv0.I a_53220_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10075 VSS word3.byte4.tinv2.I a_10020_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10076 VDD buf_in15.inv0.O buf_in15.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10077 a_20820_4840# word4.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10078 VDD word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10079 a_101600_12184# a_100810_11904# a_101430_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10080 buf_in10.inv1.O buf_in10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10081 VDD word7.byte2.tinv6.I a_124680_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10082 VSS a_149700_306# a_151260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10083 VSS a_14620_9548# a_13620_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10084 VSS buf_in6.inv0.O buf_in6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10085 a_146100_7976# word6.byte1.tinv1.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10086 a_20820_1704# word2.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10087 VDD buf_in29.inv0.O buf_in29.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10088 a_55380_11764# a_55170_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10089 a_151030_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10090 a_141060_5492# a_140850_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10091 VSS word8.byte4.tinv7.I a_28020_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10092 a_40150_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10093 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10094 VSS CLK word1.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10095 a_149700_9714# buf_out6.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10096 a_116040_2356# a_115830_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10097 VSS buf_in30.inv0.O buf_in30.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10098 Do26_buf buf_out27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10099 VSS a_55380_11764# a_55340_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10100 a_141060_2356# a_140850_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10101 a_104310_190# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10102 a_40150_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10103 buf_in21.inv1.O buf_in21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10104 word8.byte2.dff_2.O word8.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10105 a_162450_4842# word4.byte1.dff_7.CLK a_162340_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10106 VSS word2.byte3.cgate0.inv1.I word2.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10107 VDD word7.buf_sel0.O word7.byte1.nand.B VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10108 VSS a_3820_6412# a_2820_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10109 buf_sel3.inv1.O buf_sel3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10110 a_108840_11764# a_108630_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10111 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10112 word6.byte1.dff_2.O word6.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10113 VSS word2.byte4.tinv4.I a_17220_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10114 VSS a_157900_140# a_156900_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10115 a_40050_5912# buf_in24.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10116 a_57820_140# word1.byte3.cgate0.inv1.O a_58050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10117 VSS word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10118 VSS word5.byte1.cgate0.nand0.B a_134580_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10119 VSS a_60420_11112# a_61980_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10120 a_125680_7928# word6.byte2.dff_7.CLK a_125910_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10121 a_117480_306# word1.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10122 a_126800_9048# a_126010_8768# a_126630_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10123 VSS a_3820_3276# a_2820_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10124 word8.byte1.dff_0.O word8.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10125 VSS a_44580_8628# word6.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10126 VDD word1.byte1.nand.B word1.byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10127 word5.byte1.tinv7.O word5.byte1.tinv1.EN a_146100_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10128 a_7420_9548# word7.byte4.cgate0.inv1.O a_7650_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10129 word8.byte3.tinv7.O buf_out17.inv0.I a_67620_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10130 VDD a_126840_10088# a_126800_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10131 a_49620_9714# word7.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10132 VSS word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10133 a_155460_680# a_155250_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10134 VDD buf_out12.inv0.O buf_out12.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10135 a_119640_11764# a_119430_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10136 VDD word4.byte1.cgate0.nand0.B word4.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10137 a_64020_7976# buf_out18.inv0.I word6.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10138 a_54550_140# word1.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10139 a_122410_8768# word6.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10140 VSS word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10141 VDD word2.byte1.cgate0.nand0.B word2.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10142 VDD a_7420_9548# a_6420_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10143 VDD a_19380_10088# word7.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10144 VDD a_60420_4840# a_61980_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10145 a_75720_306# word1.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10146 word2.byte1.inv_and.O word2.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10147 word4.byte1.dff_3.O word4.byte1.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10148 VSS a_1380_10088# a_1340_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10149 VSS word6.byte3.tinv4.I a_56820_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10150 VSS a_106680_306# a_108240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10151 VDD a_60420_1704# a_61980_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10152 VDD buf_out32.inv0.O Do31_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10153 Do17_buf buf_out18.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10154 buf_in5.inv1.O buf_in5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10155 a_119640_8628# a_119430_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10156 VSS a_21820_11064# a_20820_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10157 a_147660_4842# a_147430_5632# a_147100_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10158 a_60420_9714# word7.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10159 a_47970_4842# a_47350_5632# a_47860_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10160 buf_we3.inv1.O buf_we3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10161 a_11580_11114# a_11350_11904# a_11020_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10162 VSS a_47020_11064# a_46020_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10163 a_113880_6578# buf_out13.inv0.I word5.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10164 a_140130_4842# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10165 a_167700_3442# word3.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10166 a_39820_140# a_40150_140# a_40050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10167 a_73020_5796# word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10168 word4.byte3.dff_5.O word4.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10169 VSS word8.byte1.cgate0.nand0.B a_73020_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10170 buf_sel4.inv1.O buf_sel4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10171 a_147660_1706# a_147430_2496# a_147100_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10172 a_115110_2776# buf_in12.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10173 VDD a_144660_6952# a_144620_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10174 a_140850_7978# word6.byte1.dff_7.CLK a_140740_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10175 a_47970_1706# a_47350_2496# a_47860_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10176 word3.byte2.tinv7.O word3.byte2.tinv6.EN a_124680_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10177 a_113880_3442# buf_out13.inv0.I word3.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10178 VDD word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10179 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10180 a_75720_7364# word5.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10181 VDD word1.byte3.buf_RE0.O word1.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10182 a_140130_1706# buf_in8.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10183 VDD buf_re.inv1.O word1.gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10184 VSS buf_sel5.inv0.O buf_sel5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10185 word2.byte3.dff_5.O word2.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10186 word7.byte2.tinv7.O buf_out15.inv0.I a_106680_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10187 VSS buf_in15.inv0.O buf_in15.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10188 a_104640_2776# word2.byte2.dff_7.CLK a_104080_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10189 VDD a_144660_3816# a_144620_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10190 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10191 a_48140_4842# word4.byte3.cgate0.inv1.O a_47970_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10192 a_158740_11114# a_156900_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10193 VDD word6.byte1.cgate0.nand0.A word6.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10194 VDD a_154300_7928# a_153300_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10195 VDD word5.byte1.cgate0.nand0.B word5.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10196 a_118710_6462# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10197 VDD word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10198 a_11860_12184# a_10020_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10199 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10200 a_75720_4228# word3.byte3.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10201 a_56820_6578# word5.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10202 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10203 a_40150_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10204 word8.byte3.cgate0.inv1.O word8.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10205 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10206 a_48140_1706# word2.byte3.cgate0.inv1.O a_47970_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10207 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.latch0.I0.O a_132960_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10208 VSS word1.byte2.tinv5.I a_121080_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10209 VDD word3.byte1.cgate0.nand0.B word3.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10210 a_115720_5912# a_113880_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10211 a_13620_6578# word5.byte4.tinv3.EN word5.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10212 a_118710_3326# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10213 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10214 word1.byte1.cgate0.inv1.I word1.byte1.cgate0.nand0.A a_134580_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10215 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10216 buf_in25.inv0.O Di24 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10217 buf_out11.inv1.O buf_out11.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10218 a_159020_12184# a_158230_11904# a_158850_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10219 a_46020_9714# buf_out23.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10220 buf_in21.inv1.O buf_in21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10221 a_7420_4792# a_7750_5632# a_7650_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10222 Do1_buf buf_out2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10223 a_154530_1090# buf_in4.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10224 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10225 a_101320_10498# a_100380_9598# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10226 VDD Di23 buf_in24.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10227 VSS word6.buf_sel0.O word6.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10228 a_112230_190# a_111610_140# a_112120_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10229 a_164100_9714# word7.byte1.tinv6.EN word7.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10230 VSS word2.byte2.cgate0.latch0.I0.O word2.byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10231 a_2820_3442# word3.byte4.tinv0.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10232 buf_sel8.inv0.I dec8.and4_7.nand1.OUT VSS VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10233 a_165660_12184# word8.byte1.dff_7.CLK a_165100_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10234 a_65020_140# a_65350_140# a_65250_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10235 VDD buf_out17.inv0.O Do16_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10236 a_125910_11114# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10237 VDD a_48180_8628# word6.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10238 a_11350_6412# word5.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10239 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10240 a_166220_190# a_165430_140# a_166050_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10241 a_147100_11064# a_147430_11904# a_147330_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10242 VSS a_146100_4840# a_147660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10243 VSS word7.byte4.buf_RE0.O word7.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10244 VDD word6.byte1.buf_RE0.I word6.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10245 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10246 a_151650_11114# a_151030_11904# a_151540_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10247 a_11350_3276# word3.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10248 a_151820_6462# a_151030_6412# a_151650_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10249 a_50850_9048# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10250 a_46020_4840# word4.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10251 a_55380_10088# a_55170_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10252 word7.byte2.dff_5.O word7.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10253 a_11250_190# buf_in29.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10254 VDD word6.gt_re3.I word6.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10255 a_112120_7362# a_110280_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10256 a_17220_9714# word7.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10257 VSS a_39820_9548# a_39720_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10258 a_110280_9714# buf_out14.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10259 VSS buf_in28.inv0.O buf_in28.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10260 a_151820_3326# a_151030_3276# a_151650_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10261 a_55060_1090# a_53220_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10262 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10263 a_46020_1704# word2.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10264 a_166260_5492# a_166050_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10265 a_112120_4226# a_110280_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10266 a_124680_11112# word8.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10267 a_122920_2776# a_121080_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10268 VSS a_48180_5492# a_48140_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10269 word7.byte2.dff_2.O word7.byte2.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10270 a_65350_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10271 a_3820_6412# word5.byte4.cgate0.inv1.O a_4050_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10272 a_40940_9598# a_40150_9548# a_40770_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10273 buf_in26.inv1.O buf_in26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10274 VSS a_151860_11764# a_151820_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10275 a_44260_190# a_42420_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10276 a_166260_2356# a_166050_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10277 buf_in20.inv1.O buf_in20.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10278 VSS CLK word6.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10279 VDD a_15780_6952# word5.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10280 word1.byte2.dff_0.O word1.byte2.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10281 VDD a_155460_680# word1.byte1.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10282 a_65350_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10283 a_134580_5796# word4.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10284 word8.byte1.tinv7.O word8.byte1.tinv2.EN a_149700_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10285 a_3820_3276# word3.byte4.cgate0.inv1.O a_4050_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10286 buf_in1.inv1.O buf_in1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10287 VSS a_51780_5492# word4.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10288 VSS a_148260_10088# a_148220_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10289 a_55380_8628# a_55170_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10290 VDD a_15780_3816# word3.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10291 VSS word4.gt_re1.O word4.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10292 VDD word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10293 a_550_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10294 VSS word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10295 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10296 a_22940_1090# word1.byte4.cgate0.inv1.O a_22770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10297 word8.byte1.nand.B word8.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10298 a_144450_7978# a_143830_8768# a_144340_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10299 VSS word5.byte2.tinv4.I a_117480_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10300 VDD word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10301 a_53220_4840# word4.byte3.tinv3.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10302 word8.byte1.tinv7.O buf_out2.inv0.I a_164100_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10303 a_119640_10088# a_119430_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10304 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10305 buf_sel1.inv0.O buf_sel1.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10306 a_15570_1706# word2.byte4.cgate0.inv1.O a_15460_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10307 a_550_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10308 VDD a_142500_6578# a_144060_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10309 a_139900_7928# a_140230_8768# a_140130_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10310 VSS word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10311 word5.byte1.nand.OUT buf_we4.inv1.O a_129540_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10312 word2.byte4.dff_7.O word2.byte4.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10313 word3.byte2.tinv7.O word3.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10314 VSS word3.byte1.cgate0.nand0.B word3.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10315 VDD buf_in11.inv0.O buf_in11.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10316 word5.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10317 VDD a_142500_3442# a_144060_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10318 VSS word5.byte1.cgate0.nand0.B word5.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10319 VSS a_153300_1704# a_154860_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10320 a_35760_7976# word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10321 a_142500_306# word1.byte1.tinv0.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10322 VSS word5.byte4.inv_and.O a_36120_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10323 VDD a_117480_306# a_119040_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10324 VDD word4.byte3.nand.OUT word4.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10325 buf_in13.inv1.O buf_in13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10326 VDD buf_out28.inv0.O Do27_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10327 a_26580_680# a_26370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10328 a_61420_9548# a_61750_9548# a_61650_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10329 VDD word2.byte3.nand.OUT word2.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10330 a_118480_6412# word5.byte2.dff_7.CLK a_118710_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10331 VSS buf_out31.inv0.O Do30_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10332 buf_in4.inv1.O buf_in4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10333 a_11580_10498# a_11350_9548# a_11020_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10334 a_155140_2776# a_153300_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10335 a_19340_6462# a_18550_6412# a_19170_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10336 VSS a_55380_2356# a_55340_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10337 VDD a_111280_6412# a_110280_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10338 a_28020_306# word1.byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10339 a_118480_3276# word3.byte2.dff_7.CLK a_118710_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10340 VSS a_26580_8628# a_26540_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10341 VDD a_54220_140# a_53220_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10342 VSS a_143500_11064# a_142500_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10343 a_19340_3326# a_18550_3276# a_19170_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10344 a_166220_5912# a_165430_5632# a_166050_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10345 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10346 VDD a_111280_3276# a_110280_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10347 a_165330_4842# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10348 a_158740_6462# a_156900_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10349 word8.byte1.cgate0.inv1.I word8.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10350 VSS a_58980_6952# a_58940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10351 a_158740_10498# a_156900_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10352 a_43420_140# word1.byte3.cgate0.inv1.O a_43650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10353 a_119320_11114# a_117480_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10354 a_111280_7928# word6.byte2.dff_7.CLK a_111510_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10355 buf_sel7.inv0.I dec8.and4_6.nand1.OUT a_75900_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10356 a_166050_7978# word6.byte1.dff_7.CLK a_165940_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10357 VDD a_8580_680# a_8540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10358 a_165330_1706# buf_in1.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10359 a_158740_3326# a_156900_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10360 a_95160_9714# word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10361 a_103080_9714# word7.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10362 VDD word4.byte2.tinv1.I a_106680_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10363 VSS buf_sel6.inv0.O buf_sel6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10364 VDD word7.byte2.cgate0.nand0.A word7.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10365 VSS a_58980_3816# a_58940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10366 a_4660_5912# a_2820_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10367 VDD word6.byte1.tinv5.I a_160500_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10368 VSS buf_in14.inv0.O buf_in14.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10369 a_40150_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10370 VSS a_116040_680# a_116000_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10371 word4.byte4.tinv7.O word4.byte4.tinv3.EN a_13620_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10372 VDD a_157900_11064# a_156900_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10373 a_64020_306# buf_out18.inv0.I word1.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10374 a_54450_7978# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10375 a_92280_12068# word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10376 VDD word2.byte2.tinv1.I a_106680_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10377 a_54450_12184# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10378 word3.byte3.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10379 VDD a_108840_5492# a_108800_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10380 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10381 word6.byte2.tinv7.O buf_out12.inv0.I a_117480_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10382 VDD word6.byte1.nand.OUT word6.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10383 a_17220_6578# word5.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10384 a_167700_306# word1.byte1.tinv7.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10385 VDD word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10386 VDD a_162660_8628# a_162620_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10387 VDD a_107680_4792# a_106680_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10388 a_151260_6462# word5.byte1.dff_7.CLK a_150700_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10389 a_119600_12184# a_118810_11904# a_119430_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10390 a_51570_6462# word5.byte3.cgate0.inv1.O a_51460_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10391 a_50950_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10392 a_4980_5492# a_4770_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10393 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10394 word5.byte3.dff_6.O word5.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10395 VDD a_108840_2356# a_108800_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10396 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10397 a_1170_190# a_550_140# a_1060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10398 a_17220_3442# word3.byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10399 VDD buf_we1.inv0.O buf_we1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10400 a_151260_3326# word3.byte1.dff_7.CLK a_150700_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10401 a_54220_11064# word8.byte3.cgate0.inv1.O a_54450_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10402 a_8540_7362# word5.byte4.cgate0.inv1.O a_8370_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10403 VDD a_107680_1656# a_106680_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10404 a_51570_3326# word3.byte3.cgate0.inv1.O a_51460_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10405 word6.byte1.tinv7.O word6.byte1.tinv6.EN a_164100_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10406 VSS word6.byte2.tinv2.I a_110280_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10407 a_167700_10500# buf_out1.inv0.I word7.byte1.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10408 word2.byte4.tinv7.O word2.byte4.tinv0.EN a_2820_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10409 VSS Di22 buf_in23.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10410 word3.byte3.dff_6.O word3.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10411 a_40380_9598# word7.byte3.cgate0.inv1.O a_39820_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10412 VDD buf_in30.inv0.O buf_in30.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10413 word8.byte3.tinv7.O word8.byte3.tinv1.EN a_46020_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10414 a_8540_4226# word3.byte4.cgate0.inv1.O a_8370_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10415 a_4150_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10416 a_125910_10498# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10417 a_4940_12184# a_4150_11904# a_4770_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10418 VSS word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10419 word1.byte1.dff_5.O word1.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10420 a_22050_7362# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10421 VDD a_166260_5492# word4.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10422 word4.byte2.dff_3.O word4.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10423 dec8.and4_0.nand0.OUT dec8.and4_6.nand0.A a_64020_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10424 VSS a_111280_7928# a_110280_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10425 VSS word2.byte1.cgate0.nand0.B word2.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10426 a_107680_11064# a_108010_11904# a_107910_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10427 a_1340_7978# word6.byte4.cgate0.inv1.O a_1170_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10428 a_19340_190# a_18550_140# a_19170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10429 VSS word1.byte3.tinv3.I a_53220_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10430 VSS a_53220_11112# a_54780_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10431 VSS a_8580_6952# word5.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10432 VDD buf_sel4.inv0.I buf_sel4.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10433 VSS CLK word8.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10434 a_112230_11114# a_111610_11904# a_112120_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10435 VDD a_107680_9548# a_106680_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10436 a_151650_9598# a_151030_9548# a_151540_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10437 a_100710_2776# buf_in16.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10438 VSS a_54220_1656# a_53220_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10439 a_1060_7362# a_120_6462# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10440 VDD a_166260_2356# word2.byte1.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10441 word1.byte2.dff_1.O word1.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10442 word2.byte2.dff_3.O word2.byte2.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10443 word3.byte2.tinv7.O word3.byte2.tinv2.EN a_110280_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10444 a_22050_4226# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10445 a_22380_1090# a_22150_140# a_21820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10446 VDD word1.byte1.cgate0.nand0.A word1.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10447 a_147430_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10448 a_144620_9048# a_143830_8768# a_144450_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10449 VSS a_8580_3816# word3.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10450 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10451 a_110280_6578# word5.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10452 a_1060_4226# a_120_3326# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10453 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10454 a_112440_11764# a_112230_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10455 a_147430_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10456 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10457 word6.byte3.buf_RE0.O word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10458 VSS a_144660_680# word1.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10459 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10460 buf_in13.inv1.O buf_in13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10461 VSS a_112440_11764# a_112400_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10462 word7.byte4.tinv7.O word7.byte4.tinv6.EN a_24420_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10463 a_28020_4840# buf_out25.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10464 word6.gt_re1.O word6.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10465 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10466 a_4770_11114# a_4150_11904# a_4660_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10467 a_140230_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10468 VSS a_11020_6412# a_10020_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10469 VDD word6.byte4.tinv7.I a_28020_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10470 a_28020_1704# buf_out25.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10471 a_450_2776# buf_in32.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10472 buf_in7.inv1.O buf_in7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10473 word1.byte2.dff_7.O word1.byte2.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10474 VSS a_11020_3276# a_10020_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10475 buf_in24.inv1.O buf_in24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10476 a_154860_190# word1.byte1.dff_7.CLK a_154300_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10477 a_118810_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10478 a_117480_4840# word4.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10479 word8.byte2.tinv7.O buf_out10.inv0.I a_124680_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10480 a_61980_7362# a_61750_6412# a_61420_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10481 VSS a_24420_7976# a_25980_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10482 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10483 word1.byte3.tinv7.O word1.byte3.tinv2.EN a_49620_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10484 a_129540_5796# word4.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10485 a_49620_11112# word8.byte3.tinv2.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10486 a_116000_7978# word6.byte2.dff_7.CLK a_115830_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10487 a_131700_7364# word5.byte1.cgate0.latch0.I0.ENB word5.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10488 VDD dec8.and4_5.nand1.B dec8.and4_1.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10489 VSS a_56820_6578# a_58380_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10490 VSS a_101640_2356# word2.byte2.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10491 word2.byte4.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10492 a_61980_4226# a_61750_3276# a_61420_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10493 VDD word1.byte1.buf_RE0.I word1.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10494 VSS word3.byte1.cgate0.nand0.B word3.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10495 a_165100_7928# a_165430_8768# a_165330_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10496 VDD a_6420_306# a_7980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10497 word3.byte1.tinv7.O word3.byte1.tinv0.EN a_142500_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10498 a_131700_4228# word3.byte1.cgate0.latch0.I0.ENB word3.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10499 a_54220_4792# word4.byte3.cgate0.inv1.O a_54450_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10500 word5.byte2.cgate0.nand0.A word5.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10501 VDD word1.gt_re3.I word1.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10502 VSS a_56820_3442# a_58380_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10503 word4.byte2.cgate0.latch0.I0.O word4.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10504 VDD buf_sel5.inv0.O buf_sel5.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10505 word8.gt_re3.I word8.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10506 VSS word3.byte4.tinv5.I a_20820_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10507 a_64020_11112# buf_out18.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10508 a_58150_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10509 a_116040_6952# a_115830_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10510 word2.byte2.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10511 a_54220_1656# word2.byte3.cgate0.inv1.O a_54450_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10512 VSS word5.byte3.cgate0.latch0.I0.O word5.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10513 word3.byte2.cgate0.nand0.A word3.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10514 a_60420_4840# buf_out19.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10515 VDD word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10516 a_40660_1090# a_39720_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10517 a_161830_8768# word6.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10518 VDD a_160500_7976# a_162060_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10519 buf_out13.inv1.O buf_out13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10520 VSS a_119640_11764# word8.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10521 buf_in27.inv0.O Di26 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10522 VSS word5.byte4.cgate0.inv1.I word5.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10523 a_116040_3816# a_115830_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10524 a_50950_5632# word4.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10525 VDD a_15780_11764# a_15740_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10526 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10527 a_60420_1704# buf_out19.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10528 Do3_buf buf_out4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10529 a_40660_11114# a_39720_11114# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10530 VDD a_141060_680# word1.byte1.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10531 a_25650_9598# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10532 a_149700_1704# word2.byte1.tinv2.EN word2.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10533 word8.byte1.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10534 a_40980_680# a_40770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10535 a_50950_2496# word2.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10536 buf_in29.inv1.O buf_in29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10537 a_36120_12068# word8.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10538 a_119320_10498# a_117480_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10539 a_118710_5912# buf_in11.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10540 word8.byte1.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10541 VDD a_20820_11112# a_22380_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10542 VSS word6.byte4.cgate0.latch0.I0.O word6.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10543 VSS word1.byte3.cgate0.nand0.A a_75360_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10544 VSS word4.byte3.buf_RE0.O word4.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10545 VDD a_111280_11064# a_110280_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10546 a_82020_5796# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10547 VSS a_121080_9714# a_122640_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10548 a_128280_9714# word7.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10549 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10550 VSS buf_ck.inv0.O CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10551 word7.gt_re0.OUT buf_sel7.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10552 a_148220_7978# word6.byte1.dff_7.CLK a_148050_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10553 word7.byte3.inv_and.O word7.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10554 word7.byte2.nand.OUT buf_we3.inv1.O a_90120_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10555 word3.gt_re3.I word3.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10556 VDD word5.byte3.dff_0.O_bar a_42420_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10557 a_35760_1092# word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10558 word8.byte2.cgate0.inv1.I word8.byte2.cgate0.nand0.A a_95160_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10559 a_144060_9048# word6.byte1.dff_7.CLK a_143500_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10560 a_150930_12184# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10561 a_44370_7978# word6.byte3.cgate0.inv1.O a_44260_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10562 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10563 a_22770_11114# word8.byte4.cgate0.inv1.O a_22660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10564 a_54220_9548# word7.byte3.cgate0.inv1.O a_54450_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10565 a_103080_9714# buf_out16.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10566 word6.byte3.dff_4.O word6.byte3.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10567 a_128280_10500# buf_out9.inv0.I word7.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10568 a_53220_3442# word3.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10569 VDD word3.byte3.dff_0.O_bar a_42420_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10570 VDD a_3820_11064# a_2820_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10571 VDD a_103080_306# a_104640_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10572 word8.byte3.dff_0.O word8.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10573 word8.byte3.dff_7.O word8.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10574 VSS a_139900_11064# a_139800_11114# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10575 word4.byte4.tinv7.O buf_out27.inv0.I a_20820_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10576 a_40980_11764# a_40770_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10577 word1.byte4.dff_3.O word1.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10578 a_140740_2776# a_139800_1706# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10579 a_11350_5632# word4.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10580 VSS a_40980_2356# a_40940_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10581 a_65580_9598# word7.byte3.cgate0.inv1.O a_65020_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10582 word2.byte4.tinv7.O buf_out27.inv0.I a_20820_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10583 VDD a_54220_9548# a_53220_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10584 a_159060_2356# a_158850_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10585 VDD Di25 buf_in26.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10586 VSS a_48180_680# a_48140_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10587 word8.byte1.tinv7.O word8.byte1.tinv7.EN a_167700_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10588 a_112230_9598# a_111610_9548# a_112120_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10589 a_115110_7362# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10590 a_58150_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10591 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10592 VSS a_112440_6952# a_112400_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10593 VSS word7.byte4.tinv1.I a_6420_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10594 a_151820_5912# a_151030_5632# a_151650_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10595 VSS buf_out3.inv0.O Do2_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10596 a_150930_4842# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10597 a_19380_5492# a_19170_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10598 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10599 a_104640_7362# a_104410_6412# a_104080_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10600 a_111510_190# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10601 VSS word2.byte3.tinv5.I a_60420_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10602 a_125910_2776# buf_in9.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10603 a_115110_4226# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10604 Do31_buf buf_out32.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10605 VDD word1.byte1.tinv5.I a_160500_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10606 VSS a_112440_3816# a_112400_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10607 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10608 a_112440_10088# a_112230_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10609 a_150930_1706# buf_in5.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10610 VSS word7.buf_ck1.I word7.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10611 a_47580_1090# a_47350_140# a_47020_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10612 a_19380_2356# a_19170_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10613 word7.byte2.cgate0.nand0.A word7.byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10614 a_550_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10615 VSS buf_we3.inv0.O buf_we3.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10616 a_104640_4226# a_104410_3276# a_104080_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10617 a_101320_9598# a_100380_9598# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10618 a_17220_1704# word2.byte4.tinv4.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10619 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10620 a_58940_4842# word4.byte3.cgate0.inv1.O a_58770_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10621 word1.byte2.tinv7.O buf_out12.inv0.I a_117480_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10622 VDD buf_sel1.inv0.O buf_sel1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10623 a_101640_680# a_101430_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10624 VDD word1.byte1.nand.OUT word1.byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10625 a_4770_9598# a_4150_9548# a_4660_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10626 VSS word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10627 a_49620_9714# word7.byte3.tinv2.EN word7.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10628 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10629 VDD word6.byte2.cgate0.nand0.A word6.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10630 word6.byte2.tinv7.O buf_out16.inv0.I a_103080_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10631 word1.byte1.cgate0.nand0.B word1.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10632 a_58940_1706# word2.byte3.cgate0.inv1.O a_58770_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10633 VSS word5.byte2.cgate0.inv1.I word5.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10634 VSS a_120_9598# a_780_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10635 a_21820_1656# a_22150_2496# a_22050_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10636 a_165430_8768# word6.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10637 buf_we4.inv0.O WE3 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X10638 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10639 VDD a_147100_6412# a_146100_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10640 VDD word7.byte4.tinv3.I a_13620_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10641 buf_in29.inv1.O buf_in29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10642 a_25420_6412# a_25750_6412# a_25650_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10643 a_51460_4842# a_49620_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10644 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10645 buf_in4.inv1.O buf_in4.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10646 a_123030_190# a_122410_140# a_122920_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10647 VDD a_147100_3276# a_146100_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10648 word6.byte2.tinv7.O word6.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10649 word1.gt_re3.I word1.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10650 a_51460_1706# a_49620_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10651 a_25420_3276# a_25750_3276# a_25650_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10652 VSS buf_in21.inv0.O buf_in21.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10653 a_162660_8628# a_162450_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10654 VDD a_151860_5492# word4.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10655 a_56820_7976# word6.byte3.tinv4.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10656 VSS a_113880_306# a_115440_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10657 a_51780_5492# a_51570_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10658 a_156900_6578# buf_out4.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10659 buf_sel3.inv0.I dec8.and4_2.nand1.OUT a_68700_13636# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10660 VSS a_126840_2356# word2.byte2.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10661 VSS word8.byte3.nand.OUT word8.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10662 VDD a_58980_8628# word6.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10663 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10664 a_20820_1704# word2.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10665 VDD a_151860_2356# word2.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10666 word7.byte3.cgate0.inv1.O word7.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10667 VSS dec8.and4_3.nand0.OUT buf_sel4.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10668 a_158130_2776# buf_in3.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10669 a_51780_2356# a_51570_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10670 word3.byte1.tinv7.O word3.byte1.tinv7.EN a_167700_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10671 a_156900_3442# buf_out4.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10672 a_58150_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10673 word5.byte1.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10674 VSS word3.byte2.tinv3.I a_113880_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10675 a_124680_4840# word4.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10676 buf_sel7.inv0.O buf_sel7.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10677 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10678 a_126840_680# a_126630_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10679 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10680 a_144340_12184# a_142500_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10681 a_19340_5912# a_18550_5632# a_19170_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10682 word5.byte1.buf_RE0.I word5.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10683 a_122920_7362# a_121080_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10684 VSS word1.byte4.buf_RE0.O word1.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10685 VDD word4.byte1.cgate0.inv1.I word4.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10686 word5.byte3.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10687 word1.gt_re1.O word1.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10688 word4.byte3.cgate0.nand0.A word4.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10689 a_18450_4842# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10690 a_154630_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10691 VDD a_15780_10088# a_15740_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10692 a_124680_1704# word2.byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10693 word7.byte4.tinv7.O word7.byte4.tinv2.EN a_10020_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10694 VSS word5.byte2.buf_RE1.I word5.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10695 buf_out12.inv1.O buf_out12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10696 VDD word1.byte4.tinv7.I a_28020_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10697 a_65860_1090# a_64020_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10698 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10699 a_40660_10498# a_39720_9598# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10700 word4.byte4.cgate0.inv1.O word4.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10701 a_119430_6462# word5.byte2.dff_7.CLK a_119320_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10702 VDD word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10703 a_158740_5912# a_156900_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10704 word2.byte3.cgate0.nand0.A word2.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10705 a_18450_1706# buf_in27.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10706 a_122920_4226# a_121080_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10707 word3.byte3.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10708 VSS a_100480_9548# a_100380_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10709 word5.byte3.tinv7.O word5.byte3.tinv4.EN a_56820_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10710 VSS a_58980_5492# a_58940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10711 VDD word6.byte4.tinv3.I a_13620_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10712 word8.gt_re3.I word8.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10713 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10714 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10715 VDD a_113880_4840# a_115440_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10716 a_119430_3326# word3.byte2.dff_7.CLK a_119320_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10717 buf_in28.inv1.O buf_in28.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10718 a_111840_12184# word8.byte2.dff_7.CLK a_111280_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10719 VDD a_20820_9714# a_22380_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10720 a_66180_680# a_65970_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10721 Do0_buf buf_out1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10722 Do22_buf buf_out23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10723 VSS a_39720_1706# a_40380_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10724 a_108240_9598# word7.byte2.dff_7.CLK a_107680_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10725 VDD a_15780_8628# a_15740_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10726 VSS a_147100_7928# a_146100_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10727 VDD a_113880_1704# a_115440_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10728 Do31_buf buf_out32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10729 VSS buf_in5.inv0.O buf_in5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10730 VSS buf_out18.inv0.O Do17_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10731 a_101600_1090# word1.byte2.dff_7.CLK a_101430_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10732 VDD a_142500_11112# a_144060_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10733 a_15570_6462# a_14950_6412# a_15460_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10734 a_155250_190# a_154630_140# a_155140_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10735 VSS a_10020_7976# a_11580_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10736 VDD a_19380_680# word1.byte4.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10737 a_90120_8932# word6.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10738 a_151260_5912# word4.byte1.dff_7.CLK a_150700_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10739 a_105030_11114# a_104410_11904# a_104920_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10740 word5.byte4.dff_7.O word5.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10741 word6.byte4.tinv7.O word6.byte4.tinv4.EN a_17220_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10742 a_51570_4842# word4.byte3.cgate0.inv1.O a_51460_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10743 VDD word4.byte4.dff_0.O_bar a_2820_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10744 VSS word2.byte1.cgate0.nand0.B a_95160_2660# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10745 a_111510_12184# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10746 a_7650_9048# buf_in30.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10747 a_64020_4840# word4.byte3.tinv6.EN word4.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10748 a_15570_3326# a_14950_3276# a_15460_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10749 word4.byte3.dff_6.O word4.byte3.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10750 VSS buf_sel1.inv0.O buf_sel1.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10751 word8.byte4.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10752 a_131700_11112# word8.byte1.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10753 word2.byte2.dff_1.O word2.byte2.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10754 VDD a_153300_6578# a_154860_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10755 VDD word2.byte4.dff_0.O_bar a_2820_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10756 word3.byte4.dff_7.O word3.byte4.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10757 VDD word5.byte3.tinv7.I a_67620_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10758 word7.byte3.dff_0.O word7.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10759 VDD a_4980_5492# a_4940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10760 word7.byte3.dff_7.O word7.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10761 word7.byte3.cgate0.inv1.I word7.byte3.cgate0.nand0.A a_73020_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10762 VDD a_153300_3442# a_154860_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10763 a_58380_4842# a_58150_5632# a_57820_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10764 a_111280_11064# word8.byte2.dff_7.CLK a_111510_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10765 VDD word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10766 word6.byte4.dff_5.O word6.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10767 word5.byte2.dff_2.O word5.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10768 word1.byte3.tinv7.O word1.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10769 VDD word3.byte3.tinv7.I a_67620_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10770 word4.byte1.nand.B word4.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10771 buf_we4.inv1.O buf_we4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10772 word7.byte1.dff_6.O word7.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10773 VSS a_10020_306# a_11580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10774 a_26540_2776# a_25750_2496# a_26370_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10775 VDD a_4980_2356# a_4940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10776 a_155140_7362# a_153300_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10777 word8.byte1.dff_6.O word8.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10778 VDD a_55380_6952# a_55340_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10779 a_58380_1706# a_58150_2496# a_57820_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10780 buf_in13.inv1.O buf_in13.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10781 word8.byte2.tinv7.O word8.byte2.tinv0.EN a_103080_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10782 word4.byte3.tinv7.O buf_out23.inv0.I a_46020_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10783 word3.byte2.dff_2.O word3.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10784 word2.byte1.nand.B word2.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10785 word8.byte2.dff_7.CLK word8.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10786 a_162660_11764# a_162450_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10787 a_119600_190# a_118810_140# a_119430_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10788 VSS a_8580_5492# word4.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10789 a_6420_7976# word6.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10790 a_155140_4226# a_153300_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10791 VSS buf_out11.inv0.O buf_out11.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10792 word7.byte4.tinv7.O word7.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10793 a_165940_2776# a_164100_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10794 VDD a_55380_3816# a_55340_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10795 VSS Di24 buf_in25.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10796 VDD a_65020_7928# a_64020_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10797 VDD a_144660_11764# word8.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10798 VDD a_150700_9548# a_149700_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10799 word2.byte3.tinv7.O buf_out23.inv0.I a_46020_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10800 VSS a_105240_8628# a_105200_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10801 VDD Di6 buf_in7.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10802 word1.byte1.dff_1.O word1.byte1.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10803 VSS word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10804 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10805 a_51460_190# a_49620_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10806 Do30_buf buf_out31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10807 a_122080_140# word1.byte2.dff_7.CLK a_122310_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10808 a_158850_190# word1.byte1.dff_7.CLK a_158740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10809 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10810 VSS a_154300_4792# a_153300_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10811 a_134580_5796# word4.byte1.cgate0.nand0.A word4.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10812 buf_in31.inv1.O buf_in31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10813 a_67620_12068# word8.byte3.tinv7.EN word8.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10814 a_113880_9714# word7.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10815 word6.byte3.tinv7.O word6.byte3.tinv2.EN a_49620_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10816 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10817 Do16_buf buf_out17.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10818 VDD word5.byte1.buf_RE0.I word5.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10819 a_65250_1090# buf_in17.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10820 word5.byte1.tinv7.O buf_out6.inv0.I a_149700_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10821 a_126520_9598# a_124680_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10822 a_22660_6462# a_20820_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10823 word4.byte2.dff_7.CLK word4.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10824 VDD buf_sel2.inv0.O buf_sel2.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10825 a_14850_11114# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10826 VDD word3.byte1.buf_RE0.I word3.byte1.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10827 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10828 word6.byte2.tinv7.O buf_out9.inv0.I a_128280_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10829 a_28020_7364# word5.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10830 a_117480_6578# word5.byte2.tinv4.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10831 word3.byte1.tinv7.O buf_out6.inv0.I a_149700_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10832 a_122640_7978# a_122410_8768# a_122080_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10833 a_22660_3326# a_20820_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10834 word6.byte3.dff_0.O word6.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10835 buf_in14.inv1.O buf_in14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10836 VDD buf_we2.inv1.O word6.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10837 a_22980_6952# a_22770_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10838 a_47020_1656# a_47350_2496# a_47250_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10839 VDD word6.byte2.nand.OUT word6.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10840 VSS word5.buf_ck1.I word5.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10841 VSS word3.byte4.nand.OUT word3.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10842 a_28020_4228# word3.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10843 a_43650_190# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10844 a_108520_1090# a_106680_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10845 a_18220_7928# a_18550_8768# a_18450_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10846 a_36120_7976# word6.byte4.cgate0.latch0.I0.ENB word6.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10847 a_149700_306# word1.byte1.tinv2.EN word1.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10848 word8.byte3.cgate0.nand0.A word8.byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10849 a_22980_3816# a_22770_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10850 VSS a_56820_4840# a_58380_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10851 a_58660_11114# a_56820_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10852 a_62540_6462# a_61750_6412# a_62370_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10853 a_19170_9598# word7.byte4.cgate0.inv1.O a_19060_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10854 a_13620_11112# word8.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10855 buf_we1.inv1.O buf_we1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10856 a_100710_7362# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10857 a_43750_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10858 word7.byte1.tinv7.O buf_out3.inv0.I a_160500_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10859 VDD word7.byte4.cgate0.inv1.I word7.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10860 a_62540_3326# a_61750_3276# a_62370_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10861 VSS buf_we2.inv0.O buf_we2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10862 a_14950_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10863 VDD a_13620_7976# a_15180_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10864 VSS a_156900_9714# a_158460_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10865 a_115210_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10866 VSS word4.byte1.buf_RE0.I word4.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10867 a_100710_4226# buf_in16.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10868 VDD buf_in18.inv0.O buf_in18.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10869 a_46020_1704# word2.byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10870 a_51740_12184# a_50950_11904# a_51570_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10871 VSS word4.gt_re3.I word4.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10872 a_73020_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10873 VSS a_7420_11064# a_6420_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10874 a_121080_11112# buf_out11.inv0.I word8.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10875 a_28020_11112# word8.byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10876 a_154300_7928# word6.byte1.dff_7.CLK a_154530_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10877 a_115210_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10878 a_112400_4842# word4.byte2.dff_7.CLK a_112230_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10879 VSS buf_sel8.inv0.O buf_sel8.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10880 a_115210_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10881 a_154630_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10882 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10883 a_146100_9714# word7.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10884 VSS word3.byte1.buf_RE1.I word3.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10885 a_8370_6462# word5.byte4.cgate0.inv1.O a_8260_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10886 VDD word4.byte1.tinv2.I a_149700_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10887 VDD word1.byte2.cgate0.nand0.A word1.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10888 word1.byte2.tinv7.O buf_out16.inv0.I a_103080_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10889 VSS word8.byte3.cgate0.inv1.I word8.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10890 a_105240_10088# a_105030_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10891 VSS word1.byte1.cgate0.nand0.B word1.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10892 a_112400_1706# word2.byte2.dff_7.CLK a_112230_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10893 a_106680_4840# buf_out15.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10894 VSS word5.byte1.buf_RE0.I word5.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10895 word4.byte2.tinv7.O word4.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10896 a_160500_7976# buf_out3.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10897 a_60420_6578# word5.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10898 VSS word7.byte4.cgate0.nand0.A a_35760_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10899 a_151030_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10900 VDD word2.byte1.tinv2.I a_149700_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10901 a_8370_3326# word3.byte4.cgate0.inv1.O a_8260_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10902 VDD a_2820_4840# a_4380_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10903 a_450_7362# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10904 VSS a_123240_680# a_123200_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10905 VSS word5.gt_re0.OUT word5.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10906 word8.byte3.dff_5.O word8.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10907 a_106680_1704# buf_out15.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X10908 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10909 buf_out16.inv1.O buf_out16.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10910 VSS a_125680_9548# a_124680_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10911 VSS a_21820_6412# a_20820_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10912 a_60420_3442# word3.byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10913 VDD word4.byte3.buf_RE0.O word4.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10914 VSS a_62580_10088# word7.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10915 VDD a_2820_1704# a_4380_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10916 a_550_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10917 a_450_4226# buf_in32.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10918 a_58980_11764# a_58770_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10919 word8.byte1.buf_RE0.I word8.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10920 Do6_buf buf_out7.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10921 a_39820_11064# a_40150_11904# a_40050_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X10922 VDD a_142500_9714# a_144060_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10923 a_780_7978# a_550_8768# a_220_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10924 VDD word2.byte3.buf_RE0.O word2.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10925 VSS a_21820_3276# a_20820_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10926 a_51570_11114# a_50950_11904# a_51460_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10927 VSS word6.byte1.tinv3.I a_153300_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10928 a_105030_9598# a_104410_9548# a_104920_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10929 VSS a_64020_1704# a_65580_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10930 VDD a_101640_6952# word5.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10931 a_58980_680# a_58770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10932 a_110280_7976# word6.byte2.tinv2.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10933 a_126800_1090# word1.byte2.dff_7.CLK a_126630_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10934 VSS buf_out22.inv0.I buf_out22.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X10935 VDD a_107680_140# a_106680_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X10936 VDD a_44580_680# word1.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10937 VDD a_101640_3816# word3.byte2.tinv0.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10938 word4.byte1.dff_4.O word4.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10939 word7.byte1.dff_7.CLK word7.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10940 a_35760_5796# word4.byte1.cgate0.nand0.B word4.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10941 a_111280_9548# word7.byte2.dff_7.CLK a_111510_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X10942 a_143730_2776# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10943 VSS word2.byte3.nand.OUT word2.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10944 word3.byte1.tinv7.O word3.byte1.tinv3.EN a_153300_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10945 a_26540_190# a_25750_140# a_26370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10946 VSS word1.byte3.tinv5.I a_60420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10947 word2.byte1.dff_4.O word2.byte1.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10948 a_101430_1706# word2.byte2.dff_7.CLK a_101320_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10949 word8.byte2.dff_6.O word8.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10950 word7.byte1.dff_6.O word7.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10951 VSS word7.byte1.buf_RE0.I word7.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10952 word1.byte2.dff_3.O word1.byte2.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X10953 a_153300_6578# word5.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10954 word6.byte3.dff_1.O word6.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10955 VDD word1.byte4.tinv3.I a_13620_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10956 VSS a_112440_5492# a_112400_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10957 VDD a_105240_11764# word8.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10958 VDD a_144660_10088# word7.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X10959 a_105030_6462# word5.byte2.dff_7.CLK a_104920_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10960 VSS a_151860_680# word1.byte1.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10961 word4.byte4.tinv7.O word4.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10962 buf_in10.inv0.O buf_in10.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10963 a_104310_9598# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X10964 buf_we1.inv1.O buf_we1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10965 a_119640_680# a_119430_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X10966 a_105030_3326# word3.byte2.dff_7.CLK a_104920_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X10967 a_119320_4842# a_117480_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10968 buf_in6.inv1.O buf_in6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10969 VSS word2.byte2.tinv1.I a_106680_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10970 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10971 word7.byte3.tinv7.O buf_out20.inv0.I a_56820_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10972 VSS word4.byte1.tinv5.I a_160500_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10973 buf_in30.inv1.O buf_in30.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10974 VSS buf_out27.inv0.I buf_out27.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X10975 a_18550_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X10976 a_140850_190# a_140230_140# a_140740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X10977 a_44260_2776# a_42420_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10978 a_119320_1706# a_117480_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10979 a_15180_12184# word8.byte4.cgate0.inv1.O a_14620_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10980 a_164100_11112# word8.byte1.tinv6.EN word8.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X10981 buf_in21.inv0.O Di20 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10982 a_14850_10498# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X10983 a_15460_9048# a_13620_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10984 VSS word6.byte3.cgate0.nand0.A a_75360_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10985 word2.byte1.cgate0.nand0.B word2.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10986 VSS word4.byte1.nand.OUT word4.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X10987 word4.byte2.tinv7.O word4.byte2.tinv4.EN a_117480_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10988 a_159020_7978# word6.byte1.dff_7.CLK a_158850_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X10989 VDD word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X10990 a_47860_6462# a_46020_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10991 VSS a_144660_2356# word2.byte1.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10992 VSS a_107680_1656# a_106680_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X10993 VDD word5.byte2.tinv5.I a_121080_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X10994 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X10995 a_44580_2356# a_44370_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X10996 word4.byte1.cgate0.nand0.B word4.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X10997 VDD EN dec8.and4_4.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X10998 a_154860_9048# word6.byte1.dff_7.CLK a_154300_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X10999 a_47860_3326# a_46020_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11000 VDD a_161500_4792# a_160500_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11001 a_43980_4842# a_43750_5632# a_43420_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11002 a_25420_4792# a_25750_5632# a_25650_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11003 VDD word7.byte2.nand.OUT word7.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11004 a_15780_8628# a_15570_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11005 VDD word3.byte2.tinv5.I a_121080_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11006 a_142500_4840# word4.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11007 a_7750_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11008 word8.byte3.tinv7.O word8.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11009 a_64020_3442# word3.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11010 a_48180_6952# a_47970_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11011 a_140740_7362# a_139800_6462# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11012 VDD word4.byte2.buf_RE1.I word4.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11013 a_92280_4840# word4.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11014 a_58660_10498# a_56820_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11015 VDD a_40980_6952# a_40940_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11016 VDD a_161500_1656# a_160500_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11017 a_43980_1706# a_43750_2496# a_43420_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11018 a_142500_1704# word2.byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11019 a_159060_6952# a_158850_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11020 a_7750_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11021 a_20820_3442# word3.byte4.tinv5.EN word3.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11022 a_26580_11764# a_26370_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11023 VDD word6.byte1.cgate0.nand0.B word6.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11024 a_1060_190# a_120_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11025 a_58150_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11026 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11027 a_55340_9048# a_54550_8768# a_55170_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11028 a_48180_3816# a_47970_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11029 VDD word2.byte2.buf_RE1.I word2.byte2.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11030 a_92280_1704# word2.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11031 a_140740_4226# a_139800_3326# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11032 VSS a_105240_10088# word7.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11033 word1.byte4.cgate0.inv1.O word1.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11034 VDD a_40980_3816# a_40940_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11035 VDD a_50620_11064# a_49620_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11036 VDD word6.byte1.buf_RE0.I word6.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11037 VDD a_50620_7928# a_49620_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11038 a_159060_3816# a_158850_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11039 a_58150_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11040 a_134580_12068# word8.byte1.cgate0.nand0.A word8.byte1.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11041 a_125910_7362# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11042 a_108010_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11043 VSS buf_in24.inv0.O buf_in24.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11044 a_151860_8628# a_151650_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11045 VSS a_106680_1704# a_108240_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11046 a_115210_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11047 word2.byte1.tinv7.O word2.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11048 a_125910_4226# buf_in9.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11049 VDD buf_in5.inv0.O buf_in5.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11050 VDD buf_out18.inv0.I buf_out18.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11051 a_119430_4842# word4.byte2.dff_7.CLK a_119320_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11052 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11053 a_149700_11112# word8.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11054 a_60420_9714# buf_out19.inv0.I word7.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11055 word8.byte4.tinv7.O buf_out29.inv0.I a_13620_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11056 a_50850_1090# buf_in21.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11057 a_28020_2660# word2.byte4.tinv7.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11058 VDD a_55380_5492# word4.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11059 word1.gt_re1.O word1.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11060 word4.gt_re1.O word4.gt_re0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11061 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11062 word1.byte2.tinv7.O buf_out9.inv0.I a_128280_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11063 a_132960_4840# word4.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11064 a_21820_6412# word5.byte4.cgate0.inv1.O a_22050_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11065 word7.byte3.dff_5.O word7.byte3.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11066 VSS word4.byte4.tinv7.I a_28020_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11067 a_155250_11114# word8.byte1.dff_7.CLK a_155140_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11068 a_103080_6578# word5.byte2.tinv0.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11069 VDD a_55380_2356# word2.byte3.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11070 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11071 VDD buf_we2.inv1.O word1.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11072 VDD word1.byte2.nand.OUT word1.byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11073 a_119040_190# word1.byte2.dff_7.CLK a_118480_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11074 a_550_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11075 VDD word5.byte1.buf_RE0.I word5.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11076 a_28020_306# word1.byte4.tinv7.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11077 a_132960_1704# word2.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11078 word3.byte1.dff_7.CLK word3.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11079 buf_out15.inv1.O buf_out15.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11080 word3.gt_re3.I word3.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11081 a_21820_3276# word3.byte4.cgate0.inv1.O a_22050_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11082 a_36120_1092# word1.byte4.cgate0.latch0.I0.ENB word1.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11083 a_42420_6578# buf_out24.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11084 a_51570_9598# a_50950_9548# a_51460_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11085 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11086 VDD word3.byte1.buf_RE0.I word3.byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11087 a_155460_11764# a_155250_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11088 VDD a_157900_6412# a_156900_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11089 a_104080_6412# a_104410_6412# a_104310_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11090 a_42420_3442# buf_out24.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11091 VDD word4.byte4.tinv2.I a_10020_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11092 VSS a_121080_11112# a_122640_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11093 VDD a_157900_3276# a_156900_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11094 VSS a_15780_11764# word8.byte4.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11095 a_104080_3276# a_104410_3276# a_104310_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11096 VDD a_126840_6952# word5.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11097 VDD word8.buf_ck1.I word8.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11098 VSS word6.byte1.cgate0.inv1.I word6.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11099 a_47250_6462# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11100 word7.byte4.dff_4.O word7.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11101 VDD word2.byte4.tinv2.I a_10020_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11102 word1.byte4.dff_5.O word1.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11103 a_158130_7362# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11104 VDD a_12180_5492# a_12140_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11105 VSS word6.gt_re3.I word6.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11106 a_100810_6412# word5.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11107 VSS a_155460_6952# a_155420_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11108 VDD buf_out2.inv0.O Do1_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11109 VSS a_55380_680# a_55340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11110 word2.byte2.cgate0.latch0.I0.O word2.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11111 VDD a_126840_3816# word3.byte2.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11112 word4.byte2.dff_2.O word4.byte2.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11113 VDD buf_out24.inv0.O Do23_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11114 a_47250_3326# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11115 word7.byte2.dff_6.O word7.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11116 a_19060_7978# a_17220_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11117 a_139900_140# word1.byte1.dff_7.CLK a_140130_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11118 word6.byte2.buf_RE1.I word6.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11119 word2.byte4.dff_0.O word2.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11120 a_158130_4226# buf_in3.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11121 a_6420_9714# word7.byte4.tinv1.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11122 VDD a_12180_2356# a_12140_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11123 VSS a_155460_3816# a_155420_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11124 a_100810_3276# word3.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11125 a_151650_4842# a_151030_5632# a_151540_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11126 a_131700_9714# word7.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11127 VDD a_119640_8628# word6.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11128 a_60420_1704# word2.byte3.tinv5.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11129 VSS word3.byte2.tinv6.I a_124680_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11130 VSS word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11131 a_158460_7978# a_158230_8768# a_157900_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11132 a_126630_1706# word2.byte2.dff_7.CLK a_126520_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11133 VDD a_105240_10088# word7.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11134 a_58770_7978# a_58150_8768# a_58660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11135 a_160500_306# buf_out3.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11136 word8.byte3.inv_and.O word8.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11137 a_144340_9598# a_142500_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11138 VSS a_44580_10088# a_44540_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11139 VSS word7.buf_ck1.I word7.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11140 word5.byte4.dff_1.O word5.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11141 a_151650_1706# a_151030_2496# a_151540_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11142 VDD word8.byte1.tinv3.I a_153300_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11143 VDD word6.byte1.cgate0.nand0.B word6.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11144 VDD word5.byte4.cgate0.nand0.A word5.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11145 a_93540_9714# word7.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11146 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11147 word6.byte1.tinv7.O buf_out7.inv0.I a_146100_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11148 word5.byte1.dff_7.CLK word5.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11149 a_8580_680# a_8370_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11150 word3.byte4.dff_1.O word3.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11151 a_8260_4842# a_6420_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11152 buf_in14.inv1.O buf_in14.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11153 VDD word3.byte4.cgate0.nand0.A word3.byte4.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11154 word5.byte1.dff_5.O word5.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11155 VDD word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11156 a_11580_2776# word2.byte4.cgate0.inv1.O a_11020_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11157 VDD a_39720_6462# a_40380_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11158 VSS a_107680_11064# a_106680_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11159 a_10020_306# word1.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11160 VSS buf_out14.inv0.O buf_out14.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11161 a_17220_9714# buf_out28.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11162 VSS a_1380_8628# a_1340_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11163 a_8260_1706# a_6420_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11164 VDD a_26580_680# a_26540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11165 word3.byte1.dff_5.O word3.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11166 a_124680_11112# word8.byte2.tinv6.EN word8.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11167 VDD a_39720_3326# a_40380_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11168 a_22660_5912# a_20820_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11169 a_8580_5492# a_8370_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11170 a_119040_9598# word7.byte2.dff_7.CLK a_118480_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11171 VSS a_157900_7928# a_156900_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11172 word8.byte2.cgate0.latch0.I0.O word8.byte2.cgate0.latch0.I0.ENB a_92280_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11173 VSS word6.byte1.buf_RE1.I word6.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11174 word7.byte1.tinv7.O buf_out5.inv0.I a_153300_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11175 VSS buf_in5.inv0.O buf_in5.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11176 word1.byte3.dff_1.O word1.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11177 a_166050_190# a_165430_140# a_165940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11178 buf_in20.inv0.O Di19 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11179 word5.byte2.dff_1.O word5.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11180 a_8580_2356# a_8370_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11181 VDD buf_in20.inv0.O buf_in20.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11182 VSS word1.byte2.nand.OUT word1.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11183 a_22980_5492# a_22770_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11184 word3.byte2.dff_1.O word3.byte2.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11185 VSS a_121080_306# a_122640_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11186 a_26540_7362# word5.byte4.cgate0.inv1.O a_26370_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11187 dec8.and4_5.nand1.OUT A2 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11188 VSS word7.gt_re1.O word7.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11189 word2.byte4.tinv7.O word2.byte4.tinv5.EN a_20820_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11190 VSS word3.byte1.tinv4.I a_156900_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11191 a_167700_4840# word4.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11192 a_62540_5912# a_61750_5632# a_62370_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11193 a_26580_10088# a_26370_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11194 a_105200_2776# a_104410_2496# a_105030_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11195 a_61650_4842# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11196 buf_sel1.inv1.O buf_sel1.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11197 a_157900_140# a_158230_140# a_158130_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11198 VSS word7.byte4.buf_RE0.O word7.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11199 word3.byte4.cgate0.nand0.A word3.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11200 a_26540_4226# word3.byte4.cgate0.inv1.O a_26370_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11201 a_140230_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11202 a_22150_9548# word7.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11203 word4.byte2.tinv7.O buf_out10.inv0.I a_124680_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11204 a_165940_7362# a_164100_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11205 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11206 word8.byte2.inv_and.O word8.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11207 a_167700_1704# word2.byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11208 a_46020_3442# word3.byte3.tinv1.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11209 a_61650_1706# buf_in18.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11210 word5.buf_sel0.O buf_sel5.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X11211 a_115210_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11212 a_108800_6462# a_108010_6412# a_108630_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11213 word1.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11214 a_165940_4226# a_164100_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11215 a_162620_9598# a_161830_9548# a_162450_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11216 VSS a_26580_6952# word5.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11217 word2.byte2.tinv7.O buf_out10.inv0.I a_124680_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11218 VSS buf_in10.inv0.O buf_in10.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11219 a_57820_11064# a_58150_11904# a_58050_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11220 VSS word5.byte3.tinv1.I a_46020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11221 VDD word4.gt_re3.I word4.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11222 a_56820_7976# word6.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11223 VSS word8.byte1.buf_RE0.I word8.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11224 a_108800_3326# a_108010_3276# a_108630_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11225 a_104920_4842# a_103080_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11226 VDD buf_in13.inv0.O buf_in13.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11227 buf_in27.inv1.O buf_in27.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11228 a_13620_7976# buf_out29.inv0.I word6.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11229 VSS a_26580_3816# word3.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11230 a_8370_4842# word4.byte4.cgate0.inv1.O a_8260_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11231 VDD word2.gt_re3.I word2.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11232 a_101600_190# a_100810_140# a_101430_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11233 VSS buf_in4.inv0.O buf_in4.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11234 a_104920_1706# a_103080_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11235 a_144620_1090# word1.byte1.dff_7.CLK a_144450_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11236 word4.byte2.tinv7.O word4.byte2.tinv0.EN a_103080_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11237 a_95160_5796# word4.byte2.cgate0.nand0.A word4.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11238 VSS a_62580_11764# a_62540_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11239 VDD a_6420_11112# a_7980_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11240 a_140850_190# word1.byte1.dff_7.CLK a_140740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11241 a_1380_10088# a_1170_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11242 a_47020_6412# word5.byte3.cgate0.inv1.O a_47250_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11243 buf_in19.inv1.O buf_in19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11244 VDD word5.byte1.buf_RE0.I word5.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11245 a_106680_6578# word5.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11246 word2.byte1.dff_2.O word2.byte1.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11247 a_150700_4792# word4.byte1.dff_7.CLK a_150930_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11248 word8.byte3.tinv7.O word8.byte3.tinv5.EN a_60420_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11249 a_2820_4840# buf_out32.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11250 word6.byte2.dff_5.O word6.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11251 word7.byte2.dff_7.CLK word7.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11252 a_125680_1656# a_126010_2496# a_125910_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11253 VSS buf_sel7.inv0.I buf_sel7.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11254 VDD word8.byte3.tinv2.I a_49620_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11255 a_116040_11764# a_115830_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11256 a_101640_6952# a_101430_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11257 VSS a_39820_7928# a_39720_7978# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11258 a_47020_3276# word3.byte3.cgate0.inv1.O a_47250_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11259 buf_in14.inv1.O buf_in14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11260 VSS a_42420_9714# a_43980_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11261 a_150700_1656# word2.byte1.dff_7.CLK a_150930_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11262 a_106680_3442# word3.byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11263 VDD word3.byte1.buf_RE0.I word3.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11264 a_67620_7364# buf_out17.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11265 VSS word5.byte1.nand.B a_78780_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11266 a_2820_1704# buf_out32.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11267 VDD word1.byte1.cgate0.nand0.B word1.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11268 VDD a_122080_9548# a_121080_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11269 a_101640_3816# a_101430_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11270 a_8370_11114# word8.byte4.cgate0.inv1.O a_8260_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11271 a_43750_6412# word5.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11272 VDD word1.byte1.buf_RE0.I word1.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11273 VDD word8.byte3.cgate0.nand0.A a_75360_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11274 a_39820_7928# word6.byte3.cgate0.inv1.O a_40050_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11275 a_40940_9048# a_40150_8768# a_40770_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11276 a_67620_4228# buf_out17.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11277 VSS a_122080_6412# a_121080_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11278 a_122410_2496# word2.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11279 a_43750_3276# word3.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11280 VDD buf_out10.inv0.O buf_out10.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11281 VDD a_24420_306# a_25980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11282 a_1380_11764# a_1170_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11283 a_126800_190# a_126010_140# a_126630_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11284 VSS a_122080_3276# a_121080_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11285 VSS a_148260_8628# a_148220_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11286 word7.byte4.cgate0.inv1.I word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11287 word6.byte4.tinv7.O word6.byte4.tinv1.EN a_6420_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11288 VSS buf_out1.inv0.O Do0_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11289 VSS buf_out23.inv0.O Do22_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11290 a_124680_1704# word2.byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11291 VDD buf_out6.inv0.I buf_out6.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11292 a_165100_140# word1.byte1.dff_7.CLK a_165330_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11293 VDD Di29 buf_in30.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11294 VDD buf_in26.inv0.O buf_in26.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11295 VSS word2.byte1.cgate0.inv1.I word2.byte1.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11296 VSS word6.byte3.buf_RE0.O word6.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11297 word6.byte1.cgate0.nand0.B word6.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11298 word2.byte3.cgate0.nand0.A word2.byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11299 a_105030_4842# word4.byte2.dff_7.CLK a_104920_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11300 VSS dec8.and4_0.nand0.OUT buf_sel1.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11301 VDD word8.byte2.tinv3.I a_113880_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11302 a_166050_190# word1.byte1.dff_7.CLK a_165940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11303 VDD a_40980_5492# word4.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11304 a_156900_9714# word7.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11305 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11306 word2.byte4.cgate0.inv1.O word2.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11307 VDD EN dec8.and4_0.nand0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11308 VDD buf_sel4.inv0.O buf_sel4.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11309 word7.byte2.tinv7.O word7.byte2.tinv3.EN a_113880_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11310 VSS word4.byte4.tinv3.I a_13620_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11311 VDD a_40980_2356# word2.byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11312 VSS a_54220_11064# a_53220_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11313 a_161830_140# word1.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11314 a_121080_306# word1.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11315 VDD word6.byte2.tinv4.I a_117480_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11316 VDD buf_sel8.inv0.I buf_sel8.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11317 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11318 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11319 a_19380_11764# a_19170_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11320 a_7980_9598# word7.byte4.cgate0.inv1.O a_7420_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11321 word6.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11322 word5.byte4.tinv7.O buf_out25.inv0.I a_28020_7364# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11323 VDD a_64020_6578# a_65580_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11324 a_61420_7928# a_61750_8768# a_61650_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11325 VSS buf_in13.inv0.O buf_in13.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11326 a_33420_9714# word7.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11327 word7.byte2.tinv7.O buf_out13.inv0.I a_113880_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11328 VDD word4.byte1.cgate0.nand0.B word4.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11329 VSS a_19380_11764# a_19340_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11330 a_165940_11114# a_164100_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11331 word6.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11332 VDD word6.byte1.cgate0.nand0.B word6.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11333 VSS word5.buf_ck1.I word5.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11334 VDD a_119640_8628# a_119600_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11335 word3.byte4.tinv7.O buf_out25.inv0.I a_28020_4228# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11336 a_162060_9598# word7.byte1.dff_7.CLK a_161500_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11337 VDD a_118480_7928# a_117480_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11338 a_50850_190# buf_in21.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11339 VSS word2.byte4.dff_0.O_bar a_2820_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11340 VDD a_64020_3442# a_65580_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11341 a_47860_5912# a_46020_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11342 VDD a_14620_4792# a_13620_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11343 a_44260_12184# a_42420_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11344 a_62370_9598# word7.byte3.cgate0.inv1.O a_62260_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11345 VDD word6.byte4.inv_and.O a_36120_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11346 VDD word2.byte1.cgate0.nand0.B word2.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11347 a_121080_7976# word6.byte2.tinv5.EN word6.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11348 a_143830_140# word1.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11349 VSS buf_out30.inv0.O Do29_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11350 a_143730_7362# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11351 VSS word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11352 VDD a_14620_1656# a_13620_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11353 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11354 VDD buf_in24.inv0.O buf_in24.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11355 VSS a_24420_11112# a_25980_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11356 VSS a_220_6412# a_120_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11357 a_101430_6462# a_100810_6412# a_101320_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11358 a_40980_680# a_40770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11359 a_48180_5492# a_47970_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11360 word6.gt_re3.I word6.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11361 a_103080_306# word1.byte2.tinv0.EN word1.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11362 a_158230_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11363 a_143730_4226# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11364 a_144060_1090# a_143830_140# a_143500_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11365 dec8.and4_7.nand1.OUT A2 a_77160_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11366 word2.byte1.nand.B word2.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11367 word6.byte4.tinv7.O word6.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11368 a_44370_190# a_43750_140# a_44260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11369 a_101430_3326# a_100810_3276# a_101320_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11370 VSS a_220_3276# a_120_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11371 a_155420_4842# word4.byte1.dff_7.CLK a_155250_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11372 word1.byte3.dff_4.O word1.byte3.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11373 VDD word1.byte1.cgate0.nand0.B word1.byte1.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11374 a_158230_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11375 word6.byte2.dff_6.O word6.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11376 word2.byte3.tinv7.O word2.byte3.tinv1.EN a_46020_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11377 a_148050_11114# word8.byte1.dff_7.CLK a_147940_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11378 a_148260_10088# a_148050_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11379 word1.byte1.tinv7.O buf_out7.inv0.I a_146100_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11380 VSS word1.byte1.tinv1.I a_146100_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11381 a_155420_1706# word2.byte1.dff_7.CLK a_155250_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11382 VSS a_48180_2356# word2.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11383 a_47350_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11384 VSS word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11385 VSS a_65020_4792# a_64020_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11386 word5.byte2.tinv7.O word5.byte2.tinv5.EN a_121080_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11387 VDD word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11388 VSS word8.gt_re1.O word8.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11389 VSS word7.byte4.tinv6.I a_24420_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11390 word8.byte3.dff_1.O word8.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11391 a_44540_7978# word6.byte3.cgate0.inv1.O a_44370_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11392 word5.byte3.tinv7.O buf_out19.inv0.I a_60420_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11393 a_154300_11064# a_154630_11904# a_154530_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11394 VSS word3.byte4.buf_RE0.O word3.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11395 VSS word5.gt_re1.O word5.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11396 word4.byte3.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11397 a_44260_7362# a_42420_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11398 a_40380_9048# word6.byte3.cgate0.inv1.O a_39820_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11399 a_4150_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11400 word3.byte3.tinv7.O buf_out19.inv0.I a_60420_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11401 VDD word8.byte1.buf_RE0.I word8.byte2.buf_RE1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11402 a_24420_9714# word7.byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11403 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11404 a_44260_4226# a_42420_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11405 VSS buf_in26.inv0.O buf_in26.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11406 VDD a_144660_6952# word5.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11407 VDD a_6420_9714# a_7980_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11408 a_153300_7976# word6.byte1.tinv3.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11409 a_44580_6952# a_44370_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11410 VDD buf_in8.inv0.O buf_in8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11411 VSS word8.byte1.cgate0.nand0.B word8.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11412 VSS word8.byte1.inv_and.O a_131700_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11413 word1.byte4.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11414 VDD buf_in29.inv0.O buf_in29.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11415 VSS word8.byte1.tinv4.I a_156900_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11416 a_66180_680# a_65970_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11417 VSS a_11020_140# a_10020_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11418 word4.byte2.tinv7.O word4.byte2.tinv7.EN a_128280_5796# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11419 a_11020_9548# a_11350_9548# a_11250_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11420 VDD a_144660_3816# word3.byte1.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11421 VSS buf_in32.inv0.O buf_in32.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11422 buf_in18.inv1.O buf_in18.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11423 a_44580_3816# a_44370_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11424 a_55380_2356# a_55170_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11425 a_78780_5796# buf_we2.inv1.O word4.byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11426 VDD a_44580_11764# word8.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11427 a_104080_4792# a_104410_5632# a_104310_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11428 VSS word4.byte2.nand.OUT word4.byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11429 VDD buf_ck.inv0.O CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11430 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11431 VSS word3.byte1.tinv0.I a_142500_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11432 a_36120_5796# word4.byte4.cgate0.latch0.I0.O word4.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11433 a_126840_6952# a_126630_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11434 a_10020_11112# buf_out30.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11435 a_144450_1706# word2.byte1.dff_7.CLK a_144340_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11436 VSS buf_ck.inv0.I buf_ck.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11437 word1.byte1.tinv7.O word1.byte1.tinv0.EN a_142500_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11438 word7.byte1.buf_RE0.I word7.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11439 VSS word3.byte2.inv_and.O a_92280_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11440 word4.byte2.tinv7.O buf_out14.inv0.I a_110280_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11441 a_47250_5912# buf_in22.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11442 word5.byte4.nand.OUT word5.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11443 VSS word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11444 word1.byte2.dff_5.O word1.byte2.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11445 a_126840_3816# a_126630_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11446 a_56820_306# word1.byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11447 VSS a_155460_5492# a_155420_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11448 a_100810_5632# word4.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11449 a_65020_7928# word6.byte3.cgate0.inv1.O a_65250_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11450 a_148050_6462# word5.byte1.dff_7.CLK a_147940_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11451 a_110280_7976# word6.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11452 word2.byte2.tinv7.O buf_out14.inv0.I a_110280_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11453 VSS buf_out16.inv0.O buf_out16.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11454 VDD word8.byte3.buf_RE0.O word8.byte3.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11455 VSS a_116040_10088# word7.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11456 word3.byte4.nand.OUT word3.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11457 VDD a_106680_6578# a_108240_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11458 VSS buf_out9.inv0.O buf_out9.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11459 a_13620_306# buf_out29.inv0.I word1.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11460 VDD buf_in9.inv0.O buf_in9.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11461 a_147330_9598# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11462 a_162660_680# a_162450_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11463 a_148050_3326# word3.byte1.dff_7.CLK a_147940_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11464 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11465 a_118810_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11466 VDD a_106680_3442# a_108240_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11467 word4.byte4.dff_1.O word4.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11468 a_61750_8768# word6.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11469 VSS word2.byte1.tinv2.I a_149700_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11470 word5.byte4.dff_3.O word5.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11471 VDD buf_out26.inv0.O Do25_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11472 VDD a_100380_7978# a_101040_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11473 VDD a_43420_6412# a_42420_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11474 a_106680_1704# word2.byte2.tinv1.EN word2.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11475 word2.byte2.tinv7.O word2.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11476 VSS a_139800_6462# a_140460_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11477 buf_in2.inv1.O buf_in2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11478 word7.byte3.tinv7.O word7.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11479 a_160500_4840# word4.byte1.tinv5.EN word4.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11480 a_67620_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11481 word3.byte4.dff_3.O word3.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11482 word4.byte1.dff_5.O word4.byte1.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11483 VSS word6.byte3.tinv6.I a_64020_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11484 VDD buf_out32.inv0.I buf_out32.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11485 VSS a_139800_3326# a_140460_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11486 VDD a_43420_3276# a_42420_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11487 VDD word5.byte1.tinv6.I a_164100_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11488 VSS word2.byte3.buf_RE0.O word2.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11489 VSS a_150700_11064# a_149700_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11490 a_19380_10088# a_19170_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11491 a_140460_11114# a_140230_11904# a_139900_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11492 VDD word7.byte1.cgate0.nand0.B word7.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11493 word1.byte1.tinv7.O word1.byte1.tinv7.EN a_167700_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11494 a_111280_1656# a_111610_2496# a_111510_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11495 a_55170_4842# a_54550_5632# a_55060_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11496 VSS word7.buf_sel0.O word7.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11497 a_58940_190# a_58150_140# a_58770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11498 word1.byte2.cgate0.latch0.I0.O word1.byte2.cgate0.latch0.I0.O a_92280_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11499 VDD word3.byte1.tinv6.I a_164100_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11500 a_126520_11114# a_124680_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11501 a_158230_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11502 a_165940_10498# a_164100_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11503 VDD a_7420_7928# a_6420_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11504 VDD word4.byte1.cgate0.nand0.B word4.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11505 word4.byte3.dff_7.O word4.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11506 buf_sel1.inv1.O buf_sel1.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11507 word8.byte4.dff_3.O word8.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11508 a_55170_1706# a_54550_2496# a_55060_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11509 a_54450_2776# buf_in20.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11510 word4.byte1.tinv7.O buf_out8.inv0.I a_142500_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11511 a_101040_190# word1.byte2.dff_7.CLK a_100480_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11512 word3.byte3.tinv7.O word3.byte3.tinv6.EN a_64020_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11513 a_10020_306# word1.byte4.tinv2.EN word1.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11514 VDD word2.byte1.cgate0.nand0.B word2.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11515 word2.byte3.dff_7.O word2.byte3.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11516 VDD a_106680_11112# a_108240_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11517 VDD word4.byte4.tinv5.I a_20820_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11518 VSS a_162660_2356# a_162620_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11519 buf_in32.inv1.O buf_in32.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11520 a_25650_9048# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11521 VSS a_148260_10088# word7.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11522 word2.byte1.tinv7.O buf_out8.inv0.I a_142500_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11523 a_61650_12184# buf_in18.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11524 VDD word6.byte3.cgate0.latch0.I0.O word6.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11525 VDD a_10020_306# a_11580_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11526 a_58050_6462# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11527 a_126800_12184# a_126010_11904# a_126630_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11528 word5.byte4.dff_0.O word5.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11529 VDD a_161500_140# a_160500_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11530 VDD word2.byte4.tinv5.I a_20820_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11531 buf_in29.inv0.O Di28 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11532 a_115440_6462# word5.byte2.dff_7.CLK a_114880_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11533 VDD a_22980_5492# a_22940_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11534 VDD word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11535 VSS word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11536 a_7650_1090# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11537 buf_re.inv0.O RE VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11538 a_53220_306# word1.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11539 VDD buf_in23.inv0.O buf_in23.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11540 a_58050_3326# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11541 a_61420_11064# word8.byte3.cgate0.inv1.O a_61650_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11542 a_126630_6462# a_126010_6412# a_126520_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11543 word3.byte4.dff_0.O word3.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11544 a_15740_9598# a_14950_9548# a_15570_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11545 VSS a_121080_7976# a_122640_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11546 a_108630_11114# word8.byte2.dff_7.CLK a_108520_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11547 VDD a_22980_2356# a_22940_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11548 a_115440_3326# word3.byte2.dff_7.CLK a_114880_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11549 VSS Di20 buf_in21.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11550 a_108800_5912# a_108010_5632# a_108630_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11551 a_126630_3326# a_126010_3276# a_126520_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11552 word8.byte3.tinv7.O word8.byte3.tinv3.EN a_53220_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11553 VSS a_123240_10088# a_123200_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11554 a_107910_4842# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11555 VSS a_26580_5492# word4.byte4.tinv7.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11556 a_161730_7978# buf_in2.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11557 a_24420_7976# word6.byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11558 VSS a_43420_7928# a_42420_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11559 a_1340_2776# a_550_2496# a_1170_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11560 a_11580_7362# a_11350_6412# a_11020_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11561 VDD word1.byte2.tinv4.I a_117480_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11562 dec8.and4_4.nand0.OUT dec8.and4_6.nand0.A a_71220_12850# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11563 VDD word7.byte3.cgate0.nand0.A word7.byte3.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11564 word2.byte4.tinv7.O word2.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11565 a_114880_11064# a_115210_11904# a_115110_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11566 a_107910_1706# buf_in14.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11567 word1.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11568 a_146100_6578# word5.byte1.tinv1.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11569 VDD a_114880_9548# a_113880_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11570 buf_sel7.inv1.O buf_sel7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11571 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11572 VSS word7.byte3.tinv2.I a_49620_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11573 a_4940_6462# a_4150_6412# a_4770_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11574 a_11580_4226# a_11350_3276# a_11020_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11575 word3.byte1.cgate0.inv1.I word3.byte1.cgate0.nand0.A a_134580_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11576 word8.byte1.dff_7.O word8.byte1.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11577 word5.byte1.buf_RE0.I word5.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11578 word5.byte2.dff_7.CLK word5.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11579 word1.buf_ck1.I CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11580 word4.gt_re3.I word4.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11581 VDD word1.byte1.cgate0.nand0.B word1.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11582 VDD a_105240_680# a_105200_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11583 a_19170_190# word1.byte4.cgate0.inv1.O a_19060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11584 VDD word1.byte4.inv_and.O a_36120_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11585 a_65580_9048# word6.byte3.cgate0.inv1.O a_65020_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11586 a_4940_3326# a_4150_3276# a_4770_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11587 a_147100_6412# a_147430_6412# a_147330_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11588 word2.gt_re3.I word2.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11589 word3.byte1.buf_RE0.I word3.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11590 VDD buf_in16.inv0.O buf_in16.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11591 VSS a_148260_11764# word8.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11592 a_53220_4840# word4.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11593 a_140230_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11594 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11595 VSS buf_in7.inv0.O buf_in7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11596 VSS a_47020_9548# a_46020_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11597 a_146100_9714# word7.byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11598 a_147100_3276# a_147430_3276# a_147330_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11599 VDD buf_out8.inv0.I buf_out8.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11600 VDD a_44580_10088# word7.byte3.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11601 a_53220_1704# word2.byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11602 a_101640_5492# a_101430_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11603 VDD buf_in28.inv0.O buf_in28.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11604 VDD buf_out1.inv0.I buf_out1.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11605 VDD a_139900_4792# a_139800_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11606 a_62260_7978# a_60420_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11607 VSS a_161500_1656# a_160500_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11608 a_142500_1704# word2.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11609 a_143830_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11610 buf_in5.inv1.O buf_in5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11611 VDD word8.byte2.tinv1.I a_106680_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11612 a_105200_7362# word5.byte2.dff_7.CLK a_105030_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11613 a_101320_9048# a_100380_7978# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11614 a_2820_6578# word5.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11615 VDD a_139900_1656# a_139800_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11616 VSS word2.byte2.buf_RE1.I word2.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11617 a_92280_2660# word2.byte2.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11618 VSS a_62580_680# a_62540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11619 a_141020_4842# word4.byte1.dff_7.CLK a_140850_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11620 VDD a_108840_5492# word4.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11621 buf_in22.inv1.O buf_in22.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11622 word1.byte3.dff_0.O word1.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11623 a_143830_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11624 VDD a_162660_8628# word6.byte1.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11625 VSS word3.byte1.tinv7.I a_167700_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11626 VSS word4.byte1.cgate0.nand0.B a_73020_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11627 a_18450_12184# buf_in27.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11628 a_105200_4226# word3.byte2.dff_7.CLK a_105030_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11629 a_131700_11112# word8.byte1.cgate0.latch0.I0.ENB word8.byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11630 word7.byte1.buf_RE0.I word7.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11631 a_62580_8628# a_62370_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11632 a_116000_2776# a_115210_2496# a_115830_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11633 a_2820_3442# word3.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11634 VDD word8.byte4.nand.OUT word8.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11635 VSS a_4980_10088# word7.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11636 a_141020_1706# word2.byte1.dff_7.CLK a_140850_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11637 VDD a_108840_2356# word2.byte2.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11638 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.latch0.I0.O a_131700_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11639 a_124680_3442# word3.byte2.tinv6.EN word3.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11640 VSS a_50620_4792# a_49620_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11641 VSS word4.byte1.buf_RE0.I word4.byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11642 VSS a_120_7978# a_780_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11643 VDD word5.byte3.inv_and.O a_75720_7364# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11644 a_18220_140# word1.byte4.cgate0.inv1.O a_18450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11645 VDD dec8.and4_5.nand1.B dec8.and4_5.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11646 word3.byte1.buf_RE1.I word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11647 word7.gt_re0.OUT buf_sel7.inv1.O a_82020_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11648 a_75360_3442# word3.byte1.cgate0.nand0.B word3.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11649 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11650 a_18220_11064# word8.byte4.cgate0.inv1.O a_18450_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11651 VDD word8.byte4.buf_RE0.O word8.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11652 a_139900_140# a_140230_140# a_140130_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11653 word3.byte1.buf_RE0.I word3.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11654 VDD word3.byte3.inv_and.O a_75720_4228# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11655 VSS word5.byte3.tinv4.I a_56820_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11656 VSS word3.byte4.cgate0.inv1.I word3.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11657 VDD word4.byte1.buf_RE0.I word4.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11658 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11659 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11660 VDD word6.byte2.cgate0.inv1.I word6.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11661 a_14950_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11662 VSS a_160500_1704# a_162060_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11663 VDD word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11664 a_65350_11904# word8.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11665 VDD word8.byte2.cgate0.inv1.I word8.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11666 a_26370_6462# word5.byte4.cgate0.inv1.O a_26260_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11667 VSS buf_out25.inv0.O Do24_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11668 buf_in10.inv1.O buf_in10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11669 a_132960_2660# word2.byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11670 VSS a_17220_11112# a_18780_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11671 VSS word8.byte1.nand.OUT word8.byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11672 VDD buf_out7.inv0.O Do6_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11673 VDD a_22980_11764# a_22940_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11674 VSS word6.byte1.buf_RE1.I word6.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11675 VDD a_124680_7976# a_126240_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11676 a_26370_3326# word3.byte4.cgate0.inv1.O a_26260_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11677 VDD a_20820_4840# a_22380_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11678 word5.byte1.dff_2.O word5.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11679 VSS a_164100_6578# a_165660_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11680 VDD a_48180_11764# a_48140_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11681 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11682 word1.byte3.dff_3.O word1.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11683 a_140460_10498# a_140230_9548# a_139900_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11684 a_125680_6412# word5.byte2.dff_7.CLK a_125910_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11685 word6.byte1.nand.B word6.buf_sel0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11686 a_15180_9598# word7.byte4.cgate0.inv1.O a_14620_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11687 VDD a_20820_1704# a_22380_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11688 word3.byte1.dff_2.O word3.byte1.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11689 a_126520_10498# a_124680_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11690 VSS a_164100_3442# a_165660_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11691 a_161500_4792# word4.byte1.dff_7.CLK a_161730_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11692 VSS word8.byte3.buf_RE0.O word8.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11693 word7.byte4.dff_3.O word7.byte4.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11694 a_125680_3276# word3.byte2.dff_7.CLK a_125910_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11695 a_112440_6952# a_112230_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11696 word6.byte1.dff_0.O word6.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11697 VSS a_53220_9714# a_54780_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11698 VSS a_66180_6952# a_66140_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11699 a_161500_1656# word2.byte1.dff_7.CLK a_161730_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11700 VSS word2.byte4.tinv2.I a_10020_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11701 VSS word7.byte3.cgate0.inv1.I word7.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11702 VDD a_106680_9714# a_108240_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11703 a_148220_2776# a_147430_2496# a_148050_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11704 a_122410_6412# word5.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11705 a_110280_306# word1.byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11706 a_112440_3816# a_112230_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11707 VSS a_100480_7928# a_100380_7978# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11708 word4.byte1.tinv7.O buf_out1.inv0.I a_167700_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11709 word6.byte1.buf_RE1.I word6.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11710 a_36120_7364# word5.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11711 VDD word4.byte2.tinv3.I a_113880_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11712 a_42420_11112# word8.byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11713 a_50620_7928# word6.byte3.cgate0.inv1.O a_50850_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11714 a_165100_140# a_165430_140# a_165330_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11715 VSS a_66180_3816# a_66140_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11716 a_42420_9714# word7.byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11717 a_4380_6462# word5.byte4.cgate0.inv1.O a_3820_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11718 VSS a_220_4792# a_120_4842# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11719 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11720 VSS buf_in14.inv0.O buf_in14.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11721 a_4150_11904# word8.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11722 a_122410_3276# word3.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11723 a_158230_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11724 word6.byte1.buf_RE0.I word6.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11725 word2.byte1.tinv7.O buf_out1.inv0.I a_167700_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11726 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11727 VDD word2.byte2.tinv3.I a_113880_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11728 a_36120_4228# word3.byte4.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11729 VSS word5.buf_sel0.O word5.byte1.nand.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11730 VDD word6.byte2.buf_RE1.I word6.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11731 a_108240_9048# word6.byte2.dff_7.CLK a_107680_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11732 a_55170_11114# word8.byte3.cgate0.inv1.O a_55060_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11733 a_61420_9548# word7.byte3.cgate0.inv1.O a_61650_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11734 a_4380_3326# word3.byte4.cgate0.inv1.O a_3820_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11735 VDD a_116040_5492# a_116000_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11736 a_75360_11112# word8.byte3.cgate0.latch0.I0.O word8.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11737 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11738 VDD word7.byte1.cgate0.inv1.I word7.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11739 a_147940_4842# a_146100_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11740 word6.byte3.tinv7.O buf_out20.inv0.I a_56820_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11741 VDD buf_in3.inv0.O buf_in3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11742 VSS word8.byte1.tinv2.I a_149700_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11743 VDD a_116040_2356# a_116000_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11744 a_13620_11112# word8.byte4.tinv3.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11745 a_147940_1706# a_146100_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11746 a_8540_190# a_7750_140# a_8370_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11747 VSS word4.byte1.cgate0.nand0.B a_134580_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11748 Do2_buf buf_out3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11749 VDD a_61420_9548# a_60420_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11750 word4.byte1.tinv7.O word4.byte1.tinv1.EN a_146100_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11751 buf_we2.inv1.O buf_we2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11752 a_49620_7976# word6.byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11753 word8.byte2.dff_0.O word8.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11754 word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.latch0.I0.ENB a_75720_10500# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11755 VSS word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11756 VSS word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11757 a_149700_6578# word5.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11758 a_28020_11112# buf_out25.inv0.I word8.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11759 a_140460_4842# a_140230_5632# a_139900_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11760 buf_we3.inv0.O WE2 VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X11761 VSS a_12180_680# word1.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11762 a_40770_4842# a_40150_5632# a_40660_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11763 word6.byte1.dff_6.O word6.byte1.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11764 a_160500_3442# word3.byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11765 VDD word5.byte2.buf_RE1.I word5.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11766 word5.byte2.tinv7.O buf_out15.inv0.I a_106680_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11767 buf_sel8.inv1.O buf_sel8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11768 word4.byte3.dff_3.O word4.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11769 a_144660_6952# a_144450_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11770 word8.byte3.cgate0.inv1.I word8.byte3.cgate0.nand0.A a_73020_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11771 a_149700_3442# word3.byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11772 word7.byte4.cgate0.inv1.O word7.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11773 a_140460_1706# a_140230_2496# a_139900_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11774 a_40770_1706# a_40150_2496# a_40660_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11775 word3.byte2.tinv7.O buf_out15.inv0.I a_106680_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11776 VDD word3.byte2.buf_RE1.I word3.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11777 VSS CLK word5.buf_ck1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11778 word2.byte3.dff_3.O word2.byte3.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11779 a_144660_3816# a_144450_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11780 word5.byte3.tinv7.O word5.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11781 VDD word1.byte3.cgate0.latch0.I0.O word1.byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11782 a_111510_6462# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11783 VDD buf_out16.inv0.I buf_out16.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X11784 a_165430_2496# word2.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11785 VDD word1.byte4.cgate0.inv1.I word1.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11786 VDD word8.gt_re3.I word8.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11787 VSS word1.gt_re1.O word1.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11788 word3.byte3.tinv7.O word3.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11789 VSS buf_out7.inv0.I buf_out7.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X11790 VSS buf_in27.inv0.O buf_in27.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11791 a_101040_6462# word5.byte2.dff_7.CLK a_100480_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11792 a_15460_1090# a_13620_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11793 a_111510_3326# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11794 a_126840_5492# a_126630_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11795 a_25750_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11796 a_167700_2660# word2.byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11797 VSS word1.byte4.buf_RE0.O word1.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11798 VDD word7.byte4.tinv5.I a_20820_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11799 a_101040_3326# word3.byte2.dff_7.CLK a_100480_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11800 VDD word7.byte3.tinv1.I a_46020_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11801 a_154860_1090# a_154630_140# a_154300_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11802 buf_in21.inv1.O buf_in21.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11803 a_126520_9048# a_124680_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11804 VDD a_48180_6952# word5.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11805 word2.byte2.tinv7.O word2.byte2.tinv6.EN a_124680_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11806 a_25750_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11807 a_148050_4842# word4.byte1.dff_7.CLK a_147940_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11808 a_15780_680# a_15570_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11809 buf_in2.inv1.O buf_in2.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11810 dec8.and4_2.nand1.OUT dec8.and4_3.nand1.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11811 a_126010_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11812 VDD a_48180_3816# word3.byte3.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11813 VSS buf_in19.inv0.O buf_in19.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11814 a_158460_11114# a_158230_11904# a_157900_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11815 a_18220_9548# word7.byte4.cgate0.inv1.O a_18450_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11816 a_155140_190# a_153300_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11817 VSS a_58980_2356# word2.byte3.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11818 a_77160_12850# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11819 VSS word2.gt_re3.I word2.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11820 word7.byte1.tinv7.O word7.byte1.tinv4.EN a_156900_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11821 a_56820_4840# word4.byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11822 VSS word7.byte2.tinv0.I a_103080_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11823 a_55340_1090# word1.byte3.cgate0.inv1.O a_55170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11824 VSS word8.gt_re3.I word8.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11825 a_123200_7978# word6.byte2.dff_7.CLK a_123030_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11826 a_13620_4840# word4.byte4.tinv3.EN word4.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11827 VSS a_143500_6412# a_142500_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11828 VDD word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11829 word4.byte4.dff_3.O word4.byte4.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11830 VDD word8.byte4.cgate0.inv1.I word8.byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11831 a_65350_9548# word7.byte3.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11832 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11833 VSS word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11834 VSS a_139800_4842# a_140460_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11835 a_117480_7976# buf_out12.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X11836 VDD word5.byte4.tinv4.I a_17220_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11837 a_108010_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11838 VSS a_143500_3276# a_142500_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11839 a_151540_12184# a_149700_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11840 VDD a_18220_9548# a_17220_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11841 a_19170_7978# word6.byte4.cgate0.inv1.O a_19060_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11842 VSS a_112440_6952# word5.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11843 VSS a_122080_140# a_121080_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11844 VDD word3.byte3.cgate0.inv1.I word3.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11845 VDD word8.byte2.buf_RE1.I word8.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11846 a_161830_11904# word8.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11847 VDD a_22980_10088# a_22940_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11848 VDD word6.buf_ck1.I word6.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11849 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11850 buf_out10.inv1.O buf_out10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11851 VDD a_48180_10088# a_48140_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11852 VDD word3.byte4.tinv4.I a_17220_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11853 VDD word4.byte4.nand.OUT word4.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11854 VSS a_112440_3816# word3.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11855 VSS a_156900_7976# a_158460_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11856 a_164100_7976# word6.byte1.tinv6.EN word6.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11857 a_55380_6952# a_55170_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11858 VDD buf_out29.inv0.O Do28_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11859 buf_in6.inv0.O Di5 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11860 a_2820_1704# word2.byte4.tinv0.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11861 VDD a_46020_4840# a_47580_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11862 VDD a_144660_11764# a_144620_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11863 VDD word2.byte4.nand.OUT word2.byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11864 buf_in26.inv1.O buf_in26.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11865 VSS a_15780_2356# a_15740_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11866 a_55380_3816# a_55170_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11867 a_144450_6462# a_143830_6412# a_144340_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11868 VDD a_46020_1704# a_47580_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11869 word6.byte3.cgate0.inv1.O word6.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11870 a_105240_8628# a_105030_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11871 Do20_buf buf_out21.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11872 VDD a_14620_140# a_13620_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X11873 VSS word6.byte4.buf_RE0.O word6.byte4.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11874 a_144450_3326# a_143830_3276# a_144340_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11875 VSS a_141060_10088# a_141020_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11876 buf_sel4.inv1.O buf_sel4.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11877 VDD a_149700_11112# a_151260_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11878 word6.byte1.dff_7.O word6.byte1.tinv7.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X11879 word5.byte1.inv_and.O word5.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11880 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11881 a_18220_140# a_18550_140# a_18450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11882 a_58050_5912# buf_in19.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11883 a_115440_5912# word4.byte2.dff_7.CLK a_114880_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11884 VSS a_62580_8628# word6.byte3.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11885 word3.byte1.inv_and.O word3.byte1.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11886 VDD word4.byte1.buf_RE1.I word4.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11887 word5.byte1.tinv7.O word5.byte1.tinv6.EN a_164100_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11888 VSS word5.byte2.tinv2.I a_110280_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11889 a_164100_11112# word8.byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11890 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11891 VSS word1.byte1.tinv3.I a_153300_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11892 a_67620_9714# word7.byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11893 VDD word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11894 a_14850_7978# buf_in28.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11895 VDD word6.byte1.buf_RE0.I word6.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11896 word2.byte4.dff_5.O word2.byte4.tinv5.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11897 VDD word2.byte1.buf_RE1.I word2.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11898 VSS a_100480_11064# a_100380_11114# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11899 a_24420_9714# word7.byte4.tinv6.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11900 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11901 VDD buf_in11.inv0.O buf_in11.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11902 VSS word5.byte3.cgate0.inv1.I word5.byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11903 word1.byte4.dff_0.O word1.byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11904 VDD word6.gt_re0.OUT word6.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11905 a_115830_9598# word7.byte2.dff_7.CLK a_115720_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11906 VDD word7.byte1.buf_RE1.I word7.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11907 a_11970_6462# word5.byte4.cgate0.inv1.O a_11860_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11908 a_58380_190# word1.byte3.cgate0.inv1.O a_57820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11909 word5.byte4.dff_6.O word5.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11910 word8.byte2.tinv7.O word8.byte2.tinv2.EN a_110280_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11911 word8.byte1.dff_7.CLK word8.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11912 VDD a_110280_7976# a_111840_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11913 a_11970_3326# word3.byte4.cgate0.inv1.O a_11860_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11914 a_36120_10500# word7.byte4.cgate0.latch0.I0.ENB word7.byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11915 word3.byte4.dff_6.O word3.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11916 a_26260_4842# a_24420_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11917 a_111280_6412# word5.byte2.dff_7.CLK a_111510_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11918 a_4940_5912# a_4150_5632# a_4770_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11919 VDD a_151860_11764# word8.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X11920 a_4050_4842# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11921 a_12140_6462# a_11350_6412# a_11970_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11922 VSS word4.byte2.tinv4.I a_117480_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11923 VDD buf_in31.inv0.O buf_in31.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11924 buf_in17.inv1.O buf_in17.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11925 VDD Di4 buf_in5.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11926 VSS word6.byte4.cgate0.inv1.I word6.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11927 a_26260_1706# a_24420_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11928 word4.byte1.nand.OUT buf_we4.inv1.O a_129540_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11929 a_111280_3276# word3.byte2.dff_7.CLK a_111510_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X11930 a_165660_4842# a_165430_5632# a_165100_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11931 a_147100_4792# a_147430_5632# a_147330_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X11932 a_4050_1706# buf_in31.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11933 a_65970_4842# a_65350_5632# a_65860_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11934 a_54450_7362# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11935 a_12140_3326# a_11350_3276# a_11970_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11936 VSS word2.byte1.cgate0.nand0.B word2.byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11937 a_151540_6462# a_149700_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11938 VSS a_51780_6952# a_51740_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11939 word4.buf_ck1.I CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11940 a_26580_5492# a_26370_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11941 word1.byte1.buf_RE1.I word1.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11942 VSS word4.byte1.cgate0.nand0.B word4.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11943 VDD buf_out20.inv0.O Do19_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11944 a_165660_1706# a_165430_2496# a_165100_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11945 VSS a_14620_1656# a_13620_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11946 VSS a_118480_4792# a_117480_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11947 VDD a_162660_6952# a_162620_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11948 a_58660_9598# a_56820_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11949 VDD a_1380_680# a_1340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11950 a_65970_1706# a_65350_2496# a_65860_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11951 a_142500_3442# word3.byte1.tinv0.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X11952 a_54450_4226# buf_in20.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11953 word4.byte1.tinv7.O buf_out5.inv0.I a_153300_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11954 VSS word4.byte4.inv_and.O a_36120_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11955 VDD word5.byte2.cgate0.latch0.I0.O word5.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11956 word1.byte1.buf_RE0.I word1.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11957 a_151540_3326# a_149700_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11958 word7.byte2.cgate0.inv1.I word7.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11959 word1.byte1.tinv7.O word1.byte1.tinv2.EN a_149700_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11960 a_26580_2356# a_26370_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11961 VSS a_51780_3816# a_51740_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X11962 VSS buf_sel6.inv0.O buf_sel6.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11963 a_104310_9048# buf_in15.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X11964 a_40940_190# a_40150_140# a_40770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11965 VSS buf_out15.inv0.I buf_out15.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X11966 a_54780_7978# a_54550_8768# a_54220_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11967 VDD word1.byte2.buf_RE1.I word1.byte2.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X11968 a_122640_2776# word2.byte2.dff_7.CLK a_122080_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X11969 VDD a_162660_3816# a_162620_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11970 a_92280_3442# word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11971 a_143830_5632# word4.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X11972 a_66140_4842# word4.byte3.cgate0.inv1.O a_65970_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11973 a_22050_11114# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11974 a_153300_7976# word6.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11975 word2.byte1.tinv7.O buf_out5.inv0.I a_153300_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11976 a_47250_11114# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X11977 VSS a_159060_10088# word7.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11978 VDD word3.byte2.cgate0.latch0.I0.O word3.byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11979 a_58980_10088# a_58770_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X11980 word1.byte3.tinv7.O buf_out20.inv0.I a_56820_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11981 VDD a_101640_5492# a_101600_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11982 a_66140_1706# word2.byte3.cgate0.inv1.O a_65970_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11983 buf_in12.inv1.O buf_in12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11984 word5.byte4.cgate0.inv1.O word5.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11985 VSS word1.byte4.cgate0.latch0.I0.O word1.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X11986 VDD a_101640_2356# a_101600_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11987 VSS a_12180_10088# word7.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X11988 VSS a_122080_11064# a_121080_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X11989 a_1340_7362# word5.byte4.cgate0.inv1.O a_1170_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11990 buf_in8.inv1.O buf_in8.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X11991 VDD word7.byte1.tinv0.I a_142500_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X11992 a_158460_10498# a_158230_9548# a_157900_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11993 a_65860_11114# a_64020_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X11994 a_95160_8932# word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11995 a_103080_7976# word6.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11996 a_108840_8628# a_108630_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X11997 a_20820_11112# word8.byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X11998 buf_in23.inv1.O buf_in23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X11999 VSS a_43420_140# a_42420_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12000 VSS a_13620_1704# a_15180_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12001 a_1340_4226# word3.byte4.cgate0.inv1.O a_1170_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12002 word1.byte3.cgate0.latch0.I0.O word1.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12003 CLK buf_ck.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12004 VDD a_46020_11112# a_47580_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12005 VSS word7.byte2.tinv7.I a_128280_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12006 word2.byte3.buf_RE0.O word2.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12007 word3.byte1.cgate0.nand0.A word3.byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12008 a_154300_1656# a_154630_2496# a_154530_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12009 a_26370_4842# word4.byte4.cgate0.inv1.O a_26260_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12010 VSS a_1380_6952# word5.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12011 VSS a_17220_6578# a_18780_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12012 a_112120_12184# a_110280_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12013 VDD a_66180_8628# word6.byte3.tinv7.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12014 a_4380_11114# a_4150_11904# a_3820_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12015 a_122410_11904# word8.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12016 a_161830_9548# word7.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12017 a_140230_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12018 VSS a_105240_8628# word6.byte2.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12019 word3.byte2.cgate0.inv1.I word3.byte2.cgate0.nand0.A a_95160_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12020 VSS a_60420_306# a_61980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12021 VSS a_17220_3442# a_18780_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12022 VSS a_1380_3816# word3.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12023 VSS a_164100_4840# a_165660_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12024 a_14620_4792# word4.byte4.cgate0.inv1.O a_14850_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12025 VSS word3.byte3.tinv3.I a_53220_3442# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12026 a_64020_4840# word4.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12027 buf_in14.inv0.O buf_in14.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12028 a_47970_11114# word8.byte3.cgate0.inv1.O a_47860_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12029 a_140230_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12030 VDD a_105240_11764# a_105200_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12031 VDD a_144660_10088# a_144620_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12032 a_14620_1656# word2.byte4.cgate0.inv1.O a_14850_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12033 VSS word5.byte4.cgate0.latch0.I0.O word5.byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12034 VSS a_57820_9548# a_56820_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12035 a_20820_4840# buf_out27.inv0.I word4.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12036 a_114880_9548# a_115210_9548# a_115110_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12037 a_64020_1704# word2.byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12038 a_112440_5492# a_112230_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12039 a_4660_12184# a_2820_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12040 VSS a_66180_5492# a_66140_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12041 a_780_2776# word2.byte4.cgate0.inv1.O a_220_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12042 a_66180_11764# a_65970_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12043 a_20820_1704# buf_out27.inv0.I word2.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12044 Do4_buf buf_out5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12045 a_108010_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12046 a_116000_7362# word5.byte2.dff_7.CLK a_115830_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12047 VDD a_149700_9714# a_151260_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12048 word1.byte2.dff_5.O word1.byte2.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12049 a_60420_306# word1.byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12050 word2.byte2.tinv7.O word2.byte2.tinv2.EN a_110280_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12051 VDD a_39820_140# a_39720_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12052 a_4380_5912# word4.byte4.cgate0.inv1.O a_3820_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12053 a_116000_4226# word3.byte2.dff_7.CLK a_115830_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12054 a_111610_9548# word7.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12055 VSS a_166260_10088# a_166220_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12056 VSS buf_out20.inv0.I buf_out20.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X12057 a_110280_4840# word4.byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12058 VSS a_148260_680# a_148220_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12059 a_108630_4842# a_108010_5632# a_108520_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12060 a_40940_1090# word1.byte3.cgate0.inv1.O a_40770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12061 a_162450_7978# a_161830_8768# a_162340_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12062 word7.byte2.cgate0.latch0.I0.O word7.byte2.cgate0.latch0.I0.O a_92280_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12063 word6.byte4.tinv7.O word6.byte4.tinv6.EN a_24420_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12064 VSS a_49620_6578# a_51180_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12065 word4.byte3.cgate0.inv1.O word4.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12066 a_4770_9598# word7.byte4.cgate0.inv1.O a_4660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12067 a_117480_306# buf_out12.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12068 VSS buf_sel1.inv0.O buf_sel1.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12069 VDD a_160500_6578# a_162060_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12070 word8.byte4.inv_and.O word8.byte4.nand.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12071 a_108630_1706# a_108010_2496# a_108520_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12072 word7.byte4.inv_and.O word7.byte4.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12073 a_40050_7978# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12074 VSS word8.byte1.cgate0.nand0.B word8.byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12075 a_103080_7976# buf_out16.inv0.I word6.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12076 VDD a_148260_680# a_148220_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12077 word2.byte3.dff_1.O word2.byte3.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12078 VSS a_49620_3442# a_51180_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12079 VDD word1.buf_ck1.I word1.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12080 word8.byte4.dff_1.O word8.byte4.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12081 VDD a_160500_3442# a_162060_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12082 word4.gt_re3.I word4.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12083 word6.byte4.dff_4.O word6.byte4.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12084 VDD word8.byte3.tinv6.I a_64020_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12085 word5.byte2.dff_4.O word5.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12086 a_13620_3442# word3.byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12087 buf_in10.inv1.O buf_in10.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12088 a_26370_190# word1.byte4.cgate0.inv1.O a_26260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12089 VDD a_151860_10088# word7.byte1.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12090 VDD a_112440_11764# word8.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12091 word2.gt_re3.I word2.gt_re1.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12092 VDD buf_in13.inv0.I buf_in13.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12093 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12094 VDD buf_in27.inv0.O buf_in27.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12095 word3.byte2.dff_4.O word3.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12096 a_15740_12184# a_14950_11904# a_15570_11114# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12097 a_132960_10500# word7.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12098 word1.byte3.cgate0.inv1.O word1.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12099 a_144660_5492# a_144450_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12100 buf_in23.inv1.O buf_in23.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12101 VSS RE buf_re.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12102 VSS Di3 buf_in4.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12103 a_25980_9598# word7.byte4.cgate0.inv1.O a_25420_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12104 word1.byte1.buf_RE0.I word1.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12105 VSS word2.byte1.cgate0.nand0.B word2.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12106 VSS a_7420_4792# a_6420_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12107 word8.byte1.inv_and.O word8.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12108 a_18550_2496# word2.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12109 a_148220_7362# word5.byte1.dff_7.CLK a_148050_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12110 word8.byte4.cgate0.latch0.I0.O word8.byte4.cgate0.latch0.I0.O a_36120_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12111 a_144340_9048# a_142500_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12112 VSS a_44580_8628# a_44540_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12113 word2.byte1.tinv7.O word2.byte1.tinv0.EN a_142500_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12114 word7.byte3.tinv7.O buf_out18.inv0.I a_64020_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12115 a_69960_12850# A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12116 a_111510_5912# buf_in13.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12117 word6.byte1.dff_3.O word6.byte1.tinv3.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12118 word5.byte4.tinv7.O buf_out32.inv0.I a_2820_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12119 VDD a_4980_11764# word8.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12120 a_22380_12184# word8.byte4.cgate0.inv1.O a_21820_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12121 VSS word2.byte4.tinv5.I a_20820_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12122 a_148220_4226# word3.byte1.dff_7.CLK a_148050_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12123 a_159020_2776# a_158230_2496# a_158850_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12124 a_61420_140# word1.byte3.cgate0.inv1.O a_61650_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12125 buf_in19.inv0.O Di18 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12126 a_22050_10498# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12127 a_47250_10498# buf_in22.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12128 a_167700_3442# word3.byte1.tinv7.EN word3.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12129 a_101040_5912# word4.byte2.dff_7.CLK a_100480_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12130 VSS word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12131 a_121080_9714# word7.byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12132 word3.byte4.tinv7.O buf_out32.inv0.I a_2820_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12133 VDD word4.byte2.tinv6.I a_124680_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12134 VSS buf_sel7.inv0.O buf_sel7.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12135 VDD word1.byte1.buf_RE0.I word1.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12136 word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B a_132960_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12137 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12138 VSS word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12139 VDD word5.byte1.cgate0.nand0.B word5.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12140 VDD word1.gt_re0.OUT word1.gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12141 a_143730_11114# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12142 a_15570_11114# a_14950_11904# a_15460_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12143 VDD word2.byte2.tinv6.I a_124680_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12144 a_10020_9714# word7.byte4.tinv2.EN word7.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12145 word5.byte2.tinv7.O word5.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12146 a_75720_3442# word3.byte3.cgate0.latch0.I0.O word3.byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12147 a_119040_9048# word6.byte2.dff_7.CLK a_118480_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12148 VDD a_126840_5492# a_126800_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12149 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12150 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12151 VDD a_125680_4792# a_124680_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12152 VDD word7.byte2.tinv0.I a_103080_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12153 VDD word3.byte1.cgate0.nand0.B word3.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12154 buf_in16.inv1.O buf_in16.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12155 a_56820_6578# word5.byte3.tinv4.EN word5.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12156 a_65860_10498# a_64020_9714# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12157 a_119600_9598# a_118810_9548# a_119430_9598# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12158 word1.byte1.inv_and.O word1.byte1.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12159 VDD a_126840_2356# a_126800_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12160 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12161 VDD a_125680_1656# a_124680_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12162 VSS word1.byte2.cgate0.inv1.I word1.byte2.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12163 VSS a_123240_680# word1.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12164 a_115720_7978# a_113880_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12165 a_11860_4842# a_10020_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12166 a_57820_6412# a_58150_6412# a_58050_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12167 VDD a_46020_9714# a_47580_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12168 a_128280_8932# word6.byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12169 a_142500_11112# word8.byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12170 a_151860_2356# a_151650_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12171 buf_in5.inv1.O buf_in5.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12172 word6.byte3.inv_and.O word6.byte3.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12173 a_11860_1706# a_10020_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12174 word6.byte2.nand.OUT buf_we3.inv1.O a_90120_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12175 word2.gt_re3.I word2.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12176 VSS buf_in22.inv0.O buf_in22.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12177 a_57820_3276# a_58150_3276# a_58050_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12178 VSS a_112440_5492# word4.byte2.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12179 a_4380_10498# a_4150_9548# a_3820_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12180 a_122410_9548# word7.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12181 a_7420_7928# word6.byte4.cgate0.inv1.O a_7650_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12182 word1.byte4.tinv7.O word1.byte4.tinv7.EN a_28020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12183 a_22150_8768# word6.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12184 a_12180_5492# a_11970_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12185 a_155460_6952# a_155250_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12186 a_54550_6412# word5.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12187 a_53220_1704# word2.byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12188 a_107680_4792# word4.byte2.dff_7.CLK a_107910_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12189 word8.byte4.tinv7.O buf_out27.inv0.I a_20820_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12190 a_156900_11112# word8.byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12191 a_40380_1090# a_40150_140# a_39820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12192 VDD a_105240_10088# a_105200_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12193 a_153300_306# word1.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12194 a_12180_2356# a_11970_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12195 a_165430_6412# word5.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12196 a_162620_9048# a_161830_8768# a_162450_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12197 a_4150_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12198 a_155460_3816# a_155250_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12199 a_73020_9714# word7.byte3.cgate0.nand0.A word7.byte3.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12200 VDD word4.byte1.tinv4.I a_156900_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12201 a_51740_4842# word4.byte3.cgate0.inv1.O a_51570_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12202 a_82020_12068# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12203 a_54550_3276# word3.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12204 VDD buf_sel8.inv0.O buf_sel8.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12205 a_107680_1656# word2.byte2.dff_7.CLK a_107910_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12206 VSS word7.gt_re3.I word7.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12207 word3.byte2.inv_and.O word3.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12208 a_162450_11114# word8.byte1.dff_7.CLK a_162340_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12209 word7.byte4.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12210 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12211 word5.byte4.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12212 a_165430_3276# word3.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12213 word4.byte4.cgate0.nand0.A word4.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12214 VDD word2.byte1.tinv4.I a_156900_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12215 a_51740_1706# word2.byte3.cgate0.inv1.O a_51570_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12216 buf_out13.inv1.O buf_out13.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12217 word7.byte3.tinv7.O word7.byte3.tinv0.EN a_42420_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12218 word3.byte4.cgate0.latch0.I0.O word3.byte4.cgate0.latch0.I0.O a_36120_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12219 a_46020_4840# buf_out23.inv0.I word4.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12220 word6.buf_sel0.O buf_sel6.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X12221 a_104410_5632# word4.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12222 VDD a_146100_7976# a_147660_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12223 a_90120_6578# word5.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12224 VDD a_159060_5492# a_159020_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12225 word2.byte4.cgate0.nand0.A word2.byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12226 word3.byte4.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12227 word8.byte2.tinv7.O word8.byte2.tinv7.EN a_128280_12068# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12228 VSS word6.byte4.tinv1.I a_6420_7976# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12229 word5.byte4.tinv7.O word5.byte4.tinv4.EN a_17220_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12230 VDD word6.byte3.tinv1.I a_46020_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12231 word8.byte1.cgate0.nand0.B word8.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12232 a_118480_140# a_118810_140# a_118710_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12233 a_46020_1704# buf_out23.inv0.I word2.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12234 word6.byte1.cgate0.latch0.I0.O word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12235 a_104410_2496# word2.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12236 VDD a_159060_2356# a_159020_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12237 buf_in29.inv1.O buf_in29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12238 a_1380_8628# a_1170_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12239 VDD a_58980_6952# word5.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12240 VSS word6.buf_ck1.I word6.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12241 VSS a_22980_11764# word8.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12242 Do23_buf buf_out24.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12243 word4.byte4.dff_2.O word4.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12244 VSS a_48180_11764# word8.byte3.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12245 VDD a_48180_8628# a_48140_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12246 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12247 VDD a_58980_3816# word3.byte3.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12248 a_19060_2776# a_17220_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12249 VSS word2.byte1.buf_RE0.I word2.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12250 VSS a_42420_7976# a_43980_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12251 a_49620_7976# word6.byte3.tinv2.EN word6.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12252 word2.byte4.dff_2.O word2.byte4.tinv2.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12253 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12254 VDD buf_out22.inv0.O Do21_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12255 a_11970_4842# word4.byte4.cgate0.inv1.O a_11860_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12256 a_149700_6578# buf_out6.inv0.I word5.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12257 VDD A1 dec8.and4_2.nand1.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12258 VDD a_51780_8628# word6.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12259 VSS a_119640_2356# word2.byte2.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12260 VSS word4.byte2.cgate0.inv1.I word4.byte2.dff_7.CLK VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12261 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12262 a_158460_2776# word2.byte1.dff_7.CLK a_157900_1656# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12263 word4.byte4.dff_6.O word4.byte4.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12264 buf_sel3.inv0.O buf_sel3.inv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12265 a_6420_6578# word5.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12266 a_58770_1706# word2.byte3.cgate0.inv1.O a_58660_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12267 VSS a_19380_680# word1.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12268 word7.byte3.cgate0.latch0.I0.O word7.byte3.cgate0.latch0.I0.O a_75720_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12269 a_53220_306# word1.byte3.tinv3.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12270 word3.byte1.tinv7.O word3.byte1.tinv5.EN a_160500_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12271 a_149700_3442# buf_out6.inv0.I word3.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12272 VDD a_14620_11064# a_13620_11112# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12273 a_118810_140# word1.byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12274 a_40050_11114# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12275 VDD a_112440_10088# word7.byte2.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12276 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12277 a_18780_4842# a_18550_5632# a_18220_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12278 word7.byte4.cgate0.inv1.I word7.byte4.cgate0.nand0.A a_33420_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12279 word6.byte3.nand.OUT word6.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12280 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12281 a_12140_5912# a_11350_5632# a_11970_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12282 VDD word8.byte1.tinv5.I a_160500_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12283 a_11250_4842# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12284 a_154530_6462# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12285 VDD a_15780_6952# a_15740_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12286 a_18780_1706# a_18550_2496# a_18220_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12287 a_100480_9548# a_100810_9548# a_100710_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12288 a_112230_6462# word5.byte2.dff_7.CLK a_112120_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12289 buf_in12.inv1.O buf_in12.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12290 a_11250_1706# buf_in29.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12291 a_151540_5912# a_149700_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12292 word5.byte3.tinv7.O word5.byte3.tinv2.EN a_49620_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12293 a_154530_3326# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12294 VSS a_51780_5492# a_51740_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12295 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12296 VSS a_114880_11064# a_113880_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12297 word1.byte2.inv_and.O word1.byte2.nand.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12298 a_104640_11114# a_104410_11904# a_104080_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12299 VDD a_15780_3816# a_15740_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12300 buf_in3.inv1.O buf_in3.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12301 a_24420_9714# buf_out26.inv0.I word7.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12302 VDD a_25420_7928# a_24420_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12303 a_112230_3326# word3.byte2.dff_7.CLK a_112120_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12304 a_143730_190# buf_in7.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12305 VDD a_4980_10088# word7.byte4.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12306 a_43650_9598# buf_in23.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12307 Do28_buf buf_out29.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12308 word2.byte1.tinv7.O word2.byte1.tinv7.EN a_167700_2660# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12309 a_36120_306# word1.byte4.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12310 VSS word2.byte2.tinv3.I a_113880_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12311 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12312 VSS a_151860_10088# a_151820_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12313 word8.byte1.tinv7.O word8.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12314 VSS Di31 buf_in32.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12315 buf_in18.inv0.O Di17 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12316 a_144060_12184# word8.byte1.dff_7.CLK a_143500_11064# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12317 word4.byte1.buf_RE0.I word4.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12318 a_104310_11114# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12319 a_143730_10498# buf_in7.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12320 a_104920_12184# a_103080_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12321 a_15570_9598# a_14950_9548# a_15460_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12322 a_7980_9048# word6.byte4.cgate0.inv1.O a_7420_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12323 word5.byte4.dff_5.O word5.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12324 VSS word7.byte1.tinv1.I a_146100_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12325 word6.byte4.tinv7.O word6.byte4.tinv2.EN a_10020_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12326 VSS word4.byte2.buf_RE1.I word4.byte2.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12327 a_220_9548# a_550_9548# a_450_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12328 a_25650_1090# buf_in25.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12329 VSS a_44580_680# word1.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12330 a_103080_306# buf_out16.inv0.I word1.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12331 a_166220_7978# word6.byte1.dff_7.CLK a_166050_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12332 a_162340_190# a_160500_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12333 a_55060_6462# a_53220_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12334 word4.byte3.tinv7.O word4.byte3.tinv4.EN a_56820_4840# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12335 buf_ck.inv0.O buf_ck.inv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12336 word3.byte4.dff_5.O word3.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12337 VDD word5.byte3.tinv5.I a_60420_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12338 a_162060_9048# word6.byte1.dff_7.CLK a_161500_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12339 a_62370_7978# word6.byte3.cgate0.inv1.O a_62260_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12340 a_55060_3326# a_53220_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12341 a_51180_4842# a_50950_5632# a_50620_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12342 a_108520_190# a_106680_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12343 a_4660_7978# a_2820_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12344 word5.byte2.dff_0.O word5.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12345 VSS a_155460_6952# word5.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12346 VSS word3.byte1.buf_RE0.I word3.byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12347 VDD word3.byte3.tinv5.I a_60420_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12348 word4.byte3.tinv7.O word4.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12349 a_17220_6578# buf_out28.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12350 VDD a_121080_306# a_122640_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12351 buf_out9.inv1.O buf_out9.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12352 a_51180_1706# a_50950_2496# a_50620_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12353 a_103080_11112# word8.byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12354 VSS a_155460_3816# word3.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12355 word3.byte2.dff_0.O word3.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12356 VDD word8.byte1.buf_RE0.I word8.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12357 VDD word6.buf_ck1.I word6.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12358 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12359 a_17220_3442# buf_out28.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12360 VSS a_17220_4840# a_18780_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12361 VSS a_1380_5492# word4.byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12362 a_65020_11064# a_65350_11904# a_65250_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12363 a_40380_190# word1.byte3.cgate0.inv1.O a_39820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12364 a_4980_8628# a_4770_7978# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12365 a_22940_6462# a_22150_6412# a_22770_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12366 buf_in25.inv1.O buf_in25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12367 VDD a_8580_11764# a_8540_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12368 a_148260_8628# a_148050_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12369 a_22940_3326# a_22150_3276# a_22770_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12370 VSS buf_in2.inv0.O buf_in2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12371 a_117480_11112# word8.byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12372 a_47350_8768# word6.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12373 word6.byte3.cgate0.inv1.I word6.byte3.cgate0.nand0.A a_73020_8932# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12374 a_122640_7362# a_122410_6412# a_122080_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12375 a_159060_680# a_158850_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12376 VDD buf_in19.inv0.O buf_in19.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12377 VSS word8.byte3.dff_0.O_bar a_42420_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12378 buf_in31.inv1.O buf_in31.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12379 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12380 a_65580_1090# a_65350_140# a_65020_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12381 word8.byte1.tinv7.O buf_out8.inv0.I a_142500_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12382 VSS a_117480_6578# a_119040_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12383 VSS Di16 buf_in17.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12384 a_122640_4226# a_122410_3276# a_122080_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12385 word7.byte2.buf_RE1.I word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12386 a_25420_140# a_25750_140# a_25650_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12387 word1.byte1.dff_7.CLK word1.byte1.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12388 VSS word5.byte1.tinv3.I a_153300_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12389 VSS a_19380_10088# a_19340_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12390 VSS a_117480_3442# a_119040_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12391 a_2820_11112# word8.byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12392 a_110280_6578# word5.byte2.tinv2.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12393 VDD word8.byte3.tinv4.I a_56820_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12394 a_123240_11764# a_123030_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12395 word6.byte2.tinv7.O buf_out11.inv0.I a_121080_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12396 a_20820_6578# word5.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12397 word7.byte3.tinv7.O word7.byte3.tinv7.EN a_67620_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12398 VSS word1.byte1.tinv5.I a_160500_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12399 buf_in12.inv1.O buf_in12.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12400 a_73020_3442# word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12401 a_39820_1656# a_40150_2496# a_40050_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12402 a_158850_9598# word7.byte1.dff_7.CLK a_158740_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12403 VDD word4.byte4.buf_RE0.O word4.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12404 VDD buf_in15.inv0.I buf_in15.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12405 VSS a_22980_10088# word7.byte4.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12406 VSS a_54220_6412# a_53220_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12407 word3.byte4.buf_RE0.O word3.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12408 a_20820_3442# word3.byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12409 VDD word6.gt_re1.O word6.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12410 VDD a_13620_6578# a_15180_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12411 a_101320_1090# a_100380_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12412 word8.gt_re1.O word8.gt_re0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12413 a_11020_7928# a_11350_8768# a_11250_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12414 a_65580_190# word1.byte3.cgate0.inv1.O a_65020_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12415 VSS word1.byte2.tinv1.I a_106680_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12416 VDD a_165100_6412# a_164100_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12417 VSS Di5 buf_in6.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12418 Do28_buf buf_out29.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12419 VSS a_49620_4840# a_51180_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12420 a_43420_6412# a_43750_6412# a_43650_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12421 VDD word2.byte4.buf_RE0.O word2.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12422 a_113880_7976# word6.byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12423 VSS a_54220_3276# a_53220_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12424 VDD a_13620_3442# a_15180_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12425 buf_in23.inv1.O buf_in23.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12426 buf_re.inv1.O buf_re.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12427 VSS a_8580_6952# a_8540_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12428 a_154300_6412# word5.byte1.dff_7.CLK a_154530_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12429 VDD a_165100_3276# a_164100_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12430 VDD a_120_190# a_780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12431 a_43420_3276# a_43750_3276# a_43650_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12432 word8.byte1.nand.OUT buf_we4.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12433 VSS buf_out21.inv0.O Do20_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12434 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12435 VSS a_8580_3816# a_8540_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12436 a_154300_3276# word3.byte1.dff_7.CLK a_154530_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12437 a_117480_4840# word4.byte2.tinv4.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12438 VSS a_149700_9714# a_151260_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12439 word4.byte2.dff_4.O word4.byte2.tinv4.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12440 a_40050_10498# buf_in24.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12441 a_44540_11114# word8.byte3.cgate0.inv1.O a_44370_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12442 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12443 VSS word4.buf_ck1.I word4.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12444 VDD word8.byte2.tinv5.I a_121080_11112# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12445 VSS dec8.and4_4.nand0.OUT buf_sel5.inv0.I VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12446 VSS word2.byte4.nand.OUT word2.byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12447 VSS a_116040_8628# word6.byte2.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12448 a_112230_190# word1.byte2.dff_7.CLK a_112120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12449 a_1170_6462# word5.byte4.cgate0.inv1.O a_1060_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12450 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12451 VDD word4.byte1.tinv0.I a_142500_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12452 VDD buf_sel7.inv0.O buf_sel7.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12453 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12454 a_147330_9048# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12455 word7.byte3.buf_RE0.O word7.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12456 VSS a_61420_11064# a_60420_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12457 VDD word5.byte1.cgate0.nand0.B word5.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12458 word1.buf_sel0.O buf_sel1.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X12459 VDD word4.byte2.inv_and.O a_92280_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12460 a_51180_11114# a_50950_11904# a_50620_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12461 a_780_7362# a_550_6412# a_220_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12462 VDD word2.byte1.tinv0.I a_142500_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12463 a_43750_11904# word8.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12464 a_104640_10498# a_104410_9548# a_104080_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12465 a_1170_3326# word3.byte4.cgate0.inv1.O a_1060_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12466 buf_in11.inv1.O buf_in11.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12467 VDD word1.byte3.tinv1.I a_46020_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12468 VDD a_144660_5492# a_144620_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12469 VDD word2.byte2.inv_and.O a_92280_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12470 VDD word3.byte1.cgate0.nand0.B word3.byte2.cgate0.inv1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12471 VSS word5.byte3.cgate0.nand0.A a_75360_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12472 a_780_4226# a_550_3276# a_220_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12473 VSS a_119640_2356# a_119600_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12474 word1.byte2.tinv7.O word1.byte2.tinv0.EN a_103080_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12475 word7.byte2.tinv7.O buf_out11.inv0.I a_121080_9714# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12476 VDD a_144660_2356# a_144620_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12477 VSS a_26580_11764# a_26540_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12478 buf_in7.inv1.O buf_in7.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12479 buf_in28.inv1.O buf_in28.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12480 word8.byte4.tinv7.O word8.byte4.tinv6.EN a_24420_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12481 a_51460_12184# a_49620_11112# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12482 a_104310_10498# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12483 a_22380_6462# word5.byte4.cgate0.inv1.O a_21820_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12484 a_126240_9598# word7.byte2.dff_7.CLK a_125680_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12485 a_146100_7976# word6.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12486 VSS a_165100_7928# a_164100_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12487 VSS word2.byte1.buf_RE1.I word2.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12488 buf_in31.inv1.O buf_in31.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12489 VDD word7.byte4.tinv1.I a_6420_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12490 VSS buf_in17.inv0.O buf_in17.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12491 VDD a_100480_140# a_100380_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12492 a_146100_306# word1.byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12493 word1.byte3.buf_RE0.O word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12494 a_22380_3326# word3.byte4.cgate0.inv1.O a_21820_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12495 VSS word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12496 VDD buf_in22.inv0.O buf_in22.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12497 word8.byte4.cgate0.inv1.O word8.byte4.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12498 word5.byte3.dff_1.O word5.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12499 VSS a_50620_140# a_49620_306# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12500 VSS word6.byte4.cgate0.nand0.A a_35760_8932# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12501 VSS word4.gt_re0.OUT word4.gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12502 VDD word7.gt_re3.I word7.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12503 VDD word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12504 VSS buf_sel2.inv0.O buf_sel2.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12505 a_118710_7978# buf_in11.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12506 word2.byte2.dff_6.O word2.byte2.tinv6.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12507 a_128280_9714# word7.byte2.tinv7.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12508 a_134580_3442# word3.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12509 word3.byte3.dff_1.O word3.byte3.tinv1.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12510 a_108240_1090# a_108010_140# a_107680_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12511 word8.byte2.tinv7.O word8.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12512 VDD word5.gt_re3.I word5.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12513 word1.byte3.nand.OUT word1.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12514 VSS a_148260_8628# word6.byte1.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12515 VDD word3.byte1.cgate0.inv1.I word3.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12516 VSS word3.gt_re1.O word3.gt_re3.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12517 a_57820_4792# a_58150_5632# a_58050_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12518 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12519 word5.byte2.dff_7.O word5.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12520 word3.byte2.dff_7.CLK word3.byte2.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12521 VDD word3.gt_re3.I word3.byte1.buf_RE0.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12522 a_44540_2776# a_43750_2496# a_44370_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12523 word8.byte2.cgate0.latch0.I0.O word8.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12524 word8.byte3.dff_3.O word8.byte3.tinv3.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12525 a_53220_3442# word3.byte3.tinv3.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12526 word4.byte3.tinv7.O buf_out18.inv0.I a_64020_4840# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12527 a_18550_6412# word5.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12528 word1.byte2.tinv7.O word1.byte2.tinv7.EN a_128280_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12529 word3.byte2.dff_7.O word3.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12530 a_15740_9048# a_14950_8768# a_15570_7978# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12531 a_155460_5492# a_155250_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12532 word8.byte2.buf_RE1.I word8.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12533 a_161500_11064# a_161830_11904# a_161730_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12534 VDD a_8580_10088# a_8540_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12535 VDD word7.byte1.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12536 a_157900_9548# a_158230_9548# a_158130_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12537 VSS buf_in10.inv0.O buf_in10.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12538 a_54550_5632# word4.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12539 buf_we1.inv0.O WE0 VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X12540 word6.byte1.dff_7.CLK word6.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12541 word2.byte3.tinv7.O buf_out18.inv0.I a_64020_1704# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12542 VSS a_123240_8628# a_123200_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12543 a_18550_3276# word3.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12544 Do24_buf buf_out25.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12545 a_112120_4842# a_110280_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12546 a_159020_7362# word5.byte1.dff_7.CLK a_158850_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12547 buf_in6.inv1.O buf_in6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12548 word1.byte1.dff_6.O word1.byte1.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12549 word2.byte1.tinv7.O word2.byte1.tinv3.EN a_153300_1704# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12550 a_115210_140# word1.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12551 VDD word7.byte1.buf_RE0.I word7.byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12552 VSS a_6420_6578# a_7980_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12553 VSS a_18220_11064# a_17220_11112# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12554 a_11350_8768# word6.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12555 VSS word6.byte1.buf_RE0.I word6.byte2.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12556 a_95160_306# word1.byte2.cgate0.nand0.A word1.byte2.cgate0.inv1.I VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12557 a_112120_1706# a_110280_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12558 a_159020_4226# word3.byte1.dff_7.CLK a_158850_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12559 a_154630_9548# word7.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12560 a_153300_4840# word4.byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12561 VSS word8.byte1.tinv6.I a_164100_11112# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12562 VSS a_6420_3442# a_7980_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12563 a_3820_4792# word4.byte4.cgate0.inv1.O a_4050_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12564 VSS word7.byte1.inv_and.O a_131700_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12565 dec8.and4_5.nand1.B A1 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12566 VDD a_15780_5492# word4.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12567 a_151820_7978# word6.byte1.dff_7.CLK a_151650_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12568 a_40660_6462# a_39720_6462# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12569 VSS a_155460_680# a_155420_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12570 VDD a_51780_11764# word8.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12571 VSS word1.byte4.tinv3.I a_13620_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12572 a_220_11064# a_550_11904# a_450_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12573 a_3820_1656# word2.byte4.cgate0.inv1.O a_4050_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12574 VDD buf_sel3.inv0.O buf_sel3.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12575 word7.byte2.cgate0.latch0.I0.O word7.byte1.cgate0.nand0.B a_93540_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12576 VSS word3.gt_re3.I word3.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12577 a_146100_7976# buf_out7.inv0.I word6.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12578 a_46020_6578# word5.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12579 VDD a_15780_2356# word2.byte4.tinv4.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12580 VSS word5.byte1.cgate0.inv1.I word5.byte1.dff_7.CLK VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12581 word7.byte2.nand.OUT buf_we3.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12582 a_40660_3326# a_39720_3326# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12583 a_11350_11904# word8.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12584 a_42420_11112# buf_out24.inv0.I word8.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12585 a_39180_9714# buf_we1.inv1.O word7.byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12586 a_550_5632# word4.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12587 VSS a_141060_6952# word5.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12588 VSS buf_in14.inv0.I buf_in14.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12589 word4.byte1.cgate0.inv1.I word4.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12590 word6.byte2.dff_7.CLK word6.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12591 a_40980_6952# a_40770_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12592 VSS word5.gt_re3.I word5.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12593 a_65020_1656# a_65350_2496# a_65250_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12594 VDD word1.buf_ck1.I word1.byte1.cgate0.nand0.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12595 a_46020_3442# word3.byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12596 a_151860_6952# a_151650_6462# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12597 word5.byte2.buf_RE1.I word5.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12598 a_126520_1090# a_124680_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12599 a_550_2496# word2.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12600 VSS a_141060_3816# word3.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12601 VDD a_142500_4840# a_144060_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12602 VSS a_220_11064# a_120_11114# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12603 word2.byte1.cgate0.inv1.I word2.byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12604 a_40980_3816# a_40770_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12605 word3.byte4.tinv7.O word3.byte4.tinv3.EN a_13620_3442# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12606 word7.byte1.buf_RE1.I word7.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12607 a_151860_3816# a_151650_3326# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12608 VDD a_142500_1704# a_144060_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12609 a_44540_10498# word7.byte3.cgate0.inv1.O a_44370_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12610 a_61750_2496# word2.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12611 word7.byte3.dff_2.O word7.byte3.tinv2.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12612 VSS a_4980_8628# word6.byte4.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12613 VSS a_100380_1706# a_101040_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12614 a_10020_9714# word7.byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12615 a_154530_5912# buf_in4.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12616 a_141020_11114# word8.byte1.dff_7.CLK a_140850_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12617 a_166220_11114# word8.byte1.dff_7.CLK a_166050_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12618 word1.byte1.dff_1.O word1.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12619 a_64020_1704# word2.byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12620 a_118480_4792# word4.byte2.dff_7.CLK a_118710_4842# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12621 a_74820_12850# EN VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12622 VDD word7.byte3.inv_and.O a_75720_10500# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12623 a_112230_4842# word4.byte2.dff_7.CLK a_112120_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12624 VDD word8.byte4.buf_RE0.O word8.byte4.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12625 VSS a_103080_6578# a_104640_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12626 a_19170_190# a_18550_140# a_19060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12627 a_51180_10498# a_50950_9548# a_50620_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12628 a_20820_1704# word2.byte4.tinv5.EN word2.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12629 a_164100_9714# word7.byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12630 word1.byte4.tinv7.O word1.byte4.tinv2.EN a_10020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12631 VDD word4.byte1.tinv7.I a_167700_4840# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12632 word1.byte2.tinv7.O buf_out11.inv0.I a_121080_306# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12633 a_123240_10088# a_123030_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12634 a_118480_1656# word2.byte2.dff_7.CLK a_118710_1706# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12635 VSS a_103080_3442# a_104640_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12636 a_124680_4840# buf_out10.inv0.I word4.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12637 VSS word5.byte1.buf_RE1.I word5.byte1.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12638 VDD a_156900_306# a_158460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12639 word7.byte3.tinv7.O word7.byte3.tinv3.EN a_53220_9714# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12640 VDD word2.byte1.tinv7.I a_167700_1704# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12641 word4.byte1.buf_RE1.I word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12642 a_165430_11904# word8.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12643 VDD word5.byte3.nand.OUT word5.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12644 a_75360_4840# word4.byte3.cgate0.latch0.I0.O word4.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12645 VDD word1.gt_re1.O word1.gt_re3.I VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12646 VDD buf_sel5.inv0.I buf_sel5.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12647 a_7650_11114# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12648 word8.byte4.dff_5.O word8.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12649 a_124680_1704# buf_out10.inv0.I word2.byte2.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12650 buf_in15.inv1.O buf_in15.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12651 a_148260_11764# a_148050_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12652 word4.byte1.buf_RE0.I word4.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12653 a_19340_7978# word6.byte4.cgate0.inv1.O a_19170_7978# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12654 VDD word6.byte3.tinv4.I a_56820_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12655 VDD word4.byte4.cgate0.inv1.I word4.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12656 word2.byte1.buf_RE1.I word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12657 word8.buf_sel0.O buf_sel8.inv1.O VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X12658 a_75360_1704# word2.byte3.cgate0.latch0.I0.O word2.byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12659 VDD word3.byte3.nand.OUT word3.byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12660 VDD a_150700_6412# a_149700_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12661 buf_in6.inv1.O buf_in6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12662 a_58770_190# word1.byte3.cgate0.inv1.O a_58660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12663 a_105240_680# a_105030_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12664 VDD a_113880_11112# a_115440_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12665 VSS a_148260_11764# a_148220_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12666 a_19060_7362# a_17220_6578# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12667 buf_in27.inv1.O buf_in27.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12668 a_15180_9048# word6.byte4.cgate0.inv1.O a_14620_7928# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12669 word2.byte1.buf_RE0.I word2.gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12670 VDD word2.byte4.cgate0.inv1.I word2.byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12671 a_158740_7978# a_156900_7976# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12672 a_55060_5912# a_53220_4840# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12673 VDD a_58980_8628# a_58940_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12674 a_47580_6462# word5.byte3.cgate0.inv1.O a_47020_6412# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12675 VDD a_150700_3276# a_149700_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12676 VDD a_119640_6952# word5.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12677 a_100480_140# a_100810_140# a_100710_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12678 a_19060_4226# a_17220_3442# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12679 a_158460_7362# a_158230_6412# a_157900_6412# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12680 a_58770_6462# a_58150_6412# a_58660_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12681 VSS buf_in21.inv0.O buf_in21.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12682 VDD a_125680_140# a_124680_306# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12683 VSS a_53220_7976# a_54780_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12684 VDD a_62580_680# word1.byte3.tinv6.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12685 a_47580_3326# word3.byte3.cgate0.inv1.O a_47020_3276# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12686 a_103080_4840# word4.byte2.tinv0.EN word4.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12687 VDD buf_in21.inv0.O buf_in21.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12688 a_6420_11112# word8.byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12689 VDD a_119640_3816# word3.byte2.tinv5.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12690 VSS a_155460_5492# word4.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12691 word4.byte2.dff_0.O word4.byte2.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12692 buf_in2.inv0.O Di1 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12693 a_8540_4842# word4.byte4.cgate0.inv1.O a_8370_4842# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12694 a_158460_4226# a_158230_3276# a_157900_3276# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12695 a_115830_11114# word8.byte2.dff_7.CLK a_115720_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12696 word2.gt_re3.I word2.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12697 a_58770_3326# a_58150_3276# a_58660_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12698 VDD word8.byte1.cgate0.inv1.I word8.byte1.dff_7.CLK VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12699 word7.byte1.nand.B word7.buf_sel0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12700 VSS Di18 buf_in19.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12701 VDD word5.byte2.tinv1.I a_106680_6578# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12702 VSS word1.byte4.cgate0.nand0.A a_35760_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12703 a_161730_2776# buf_in2.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12704 a_8540_1706# word2.byte4.cgate0.inv1.O a_8370_1706# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12705 word8.byte1.buf_RE0.I word8.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12706 a_151260_7978# a_151030_8768# a_150700_7928# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12707 a_51570_7978# a_50950_8768# a_51460_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12708 a_117480_3442# word3.byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12709 VDD word3.byte2.tinv1.I a_106680_3442# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12710 a_22940_5912# a_22150_5632# a_22770_4842# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12711 word7.byte1.cgate0.nand0.B word7.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12712 a_22050_4842# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12713 word8.byte4.cgate0.inv1.I word8.byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12714 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12715 word6.byte3.dff_6.O word6.byte3.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12716 a_129540_3442# word3.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12717 a_122080_11064# a_122410_11904# a_122310_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12718 a_220_140# a_550_140# a_450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12719 a_22150_140# word1.byte4.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12720 VSS word1.byte3.nand.OUT word1.byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12721 a_123030_6462# word5.byte2.dff_7.CLK a_122920_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12722 a_22050_1706# buf_in26.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12723 a_1060_4842# a_120_4842# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12724 word3.byte1.cgate0.nand0.B word3.buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12725 word6.byte1.tinv7.O word6.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12726 a_147430_5632# word4.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12727 a_122310_9598# buf_in10.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12728 VDD word6.buf_sel0.O word6.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12729 a_1060_1706# a_120_1706# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12730 a_123030_3326# word3.byte2.dff_7.CLK a_122920_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12731 a_147430_2496# word2.byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12732 a_6420_7976# word6.byte4.tinv1.EN word6.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12733 VSS a_117480_4840# a_119040_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12734 Do5_buf buf_out6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12735 VSS a_155460_11764# word8.byte1.tinv4.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12736 a_111840_9598# word7.byte2.dff_7.CLK a_111280_9548# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12737 a_92280_11112# word8.byte2.inv_and.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12738 a_131700_8932# word6.byte1.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12739 VSS a_150700_7928# a_149700_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12740 VSS word2.byte2.tinv6.I a_124680_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12741 a_153300_9714# word7.byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12742 VDD a_8580_8628# word6.byte4.tinv2.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12743 VSS buf_in5.inv0.O buf_in5.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12744 VSS buf_in26.inv0.O buf_in26.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12745 a_62260_2776# a_60420_1704# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12746 VDD a_51780_10088# word7.byte3.tinv3.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12747 VSS word6.buf_ck1.I word6.byte1.cgate0.nand0.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12748 word8.byte4.buf_RE0.O word8.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12749 VDD a_18220_6412# a_17220_6578# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12750 a_104310_1090# buf_in15.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12751 a_93540_8932# word6.byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12752 word2.byte1.buf_RE0.I word2.gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12753 word4.byte1.dff_7.CLK word4.byte1.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12754 VDD word8.byte1.buf_RE1.I word8.byte1.tinv7.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12755 a_65860_6462# a_64020_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12756 VSS a_162660_2356# word2.byte1.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12757 VSS a_125680_1656# a_124680_1704# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12758 a_11350_9548# word7.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12759 a_113880_9714# word7.byte2.tinv3.EN word7.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12760 a_62580_2356# a_62370_1706# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12761 VDD a_18220_3276# a_17220_3442# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12762 word5.byte1.tinv7.O word5.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12763 a_25650_12184# buf_in25.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12764 a_65860_3326# a_64020_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12765 a_61980_4842# a_61750_5632# a_61420_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12766 a_43420_4792# a_43750_5632# a_43650_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12767 buf_sel5.inv1.O buf_sel5.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12768 a_43980_11114# a_43750_11904# a_43420_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12769 a_160500_4840# word4.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12770 word5.byte4.tinv7.O word5.byte4.tinv1.EN a_6420_6578# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12771 VSS a_8580_5492# a_8540_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12772 a_75720_9714# word7.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12773 a_60420_306# word1.byte3.tinv5.EN word1.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12774 VSS word1.buf_sel0.O word1.byte1.nand.B VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12775 VSS word3.byte3.buf_RE0.O word3.byte3.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12776 a_47350_140# word1.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12777 word3.byte1.tinv7.O word3.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12778 a_82020_3442# buf_re.inv1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12779 VSS a_154300_9548# a_153300_9714# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12780 a_28020_7364# buf_out25.inv0.I word5.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12781 a_66180_6952# a_65970_6462# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12782 a_90120_12068# word8.byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12783 a_61980_1706# a_61750_2496# a_61420_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12784 VSS word7.byte1.cgate0.nand0.B a_33420_9714# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12785 a_160500_1704# word2.byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12786 VSS word5.byte3.buf_RE0.O word5.byte3.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12787 a_25420_11064# word8.byte4.cgate0.inv1.O a_25650_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12788 VDD CLK word6.buf_ck1.I VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12789 word5.byte1.cgate0.nand0.B word5.buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12790 VDD buf_we2.inv1.O word8.byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12791 a_143500_9548# a_143830_9548# a_143730_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12792 a_101600_6462# a_100810_6412# a_101430_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12793 a_66180_3816# a_65970_3326# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12794 a_28020_4228# buf_out25.inv0.I word3.byte4.tinv7.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12795 a_155250_6462# word5.byte1.dff_7.CLK a_155140_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12796 VSS a_19380_6952# word5.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12797 VSS a_123240_10088# word7.byte2.tinv6.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12798 word8.byte4.tinv7.O word8.byte4.tinv4.EN a_17220_11112# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12799 a_101600_11114# word8.byte2.dff_7.CLK a_101430_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12800 a_141020_10498# word7.byte1.dff_7.CLK a_140850_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12801 a_155250_3326# word3.byte1.dff_7.CLK a_155140_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12802 a_101600_3326# a_100810_3276# a_101430_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12803 a_166220_10498# word7.byte1.dff_7.CLK a_166050_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12804 VSS a_19380_3816# word3.byte4.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12805 a_126010_8768# word6.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12806 a_116040_5492# a_115830_4842# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12807 a_1170_4842# word4.byte4.cgate0.inv1.O a_1060_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12808 VSS buf_out24.inv0.O Do23_buf VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12809 VDD a_56820_7976# a_58380_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12810 VSS a_124680_1704# a_126240_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12811 VSS word6.gt_re1.O word6.gt_re3.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12812 a_150930_190# buf_in5.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12813 VSS word2.byte1.tinv4.I a_156900_1704# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12814 VDD buf_out5.inv0.O Do4_buf VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12815 VDD buf_in17.inv0.O buf_in17.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12816 a_116040_2356# a_115830_1706# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12817 VSS word6.byte4.buf_RE0.O word6.byte4.tinv7.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12818 VDD a_105240_680# word1.byte2.tinv1.I VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X12819 word2.byte4.cgate0.nand0.A word2.byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12820 VDD a_55380_11764# a_55340_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12821 word4.byte1.tinv7.O word4.byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12822 a_46020_1704# word2.byte3.tinv1.EN word2.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12823 a_100810_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12824 word4.buf_sel0.O buf_sel4.inv1.O VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X12825 a_126010_11904# word8.byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12826 a_141060_680# a_140850_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12827 a_146100_306# buf_out7.inv0.I word1.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12828 buf_in19.inv1.O buf_in19.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12829 a_75720_12068# word8.byte3.inv_and.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12830 a_7650_10498# buf_in30.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12831 VSS a_18220_7928# a_17220_7976# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12832 a_39820_6412# word5.byte3.cgate0.inv1.O a_40050_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12833 word5.byte2.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12834 word2.byte1.dff_0.O word2.byte1.tinv0.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12835 word7.byte4.dff_5.O word7.byte4.tinv5.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12836 a_108840_11764# a_108630_11114# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12837 a_148260_10088# a_148050_9598# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X12838 VSS word1.byte3.cgate0.inv1.I word1.byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12839 VSS word4.byte3.tinv1.I a_46020_4840# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12840 VDD word7.byte1.buf_RE0.I word7.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12841 a_121080_6578# word5.byte2.tinv5.EN word5.byte2.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12842 VSS a_51780_680# word1.byte3.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12843 word1.byte2.dff_7.CLK word1.byte2.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12844 buf_sel6.inv1.O buf_sel6.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12845 VSS word1.gt_re3.I word1.byte1.buf_RE0.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12846 VDD a_60420_11112# a_61980_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12847 buf_in14.inv1.O buf_in14.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12848 word3.byte2.cgate0.latch0.I0.O word3.byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12849 a_39820_3276# word3.byte3.cgate0.inv1.O a_40050_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12850 a_22380_5912# word4.byte4.cgate0.inv1.O a_21820_4792# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12851 VSS word5.byte1.cgate0.latch0.I0.O word5.byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12852 buf_sel6.inv1.O buf_sel6.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12853 VDD a_113880_9714# a_115440_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12854 word5.byte3.cgate0.inv1.O word5.byte3.cgate0.inv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12855 a_50620_1656# a_50950_2496# a_50850_2776# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12856 word8.byte1.dff_0.O word8.byte1.tinv0.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12857 a_60420_6578# buf_out19.inv0.I word5.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12858 word3.byte4.tinv7.O word3.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12859 word5.byte1.dff_1.O word5.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12860 word5.gt_re3.I word5.gt_re1.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12861 VDD word4.byte1.buf_RE0.I word4.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12862 a_115720_190# a_113880_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12863 a_122080_6412# a_122410_6412# a_122310_6462# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12864 VSS buf_in12.inv0.O buf_in12.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12865 word5.byte4.tinv7.O word5.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12866 a_60420_3442# buf_out19.inv0.I word3.byte3.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12867 word3.byte1.dff_1.O word3.byte1.tinv1.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12868 VDD word2.byte1.buf_RE0.I word2.byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12869 buf_in8.inv1.O buf_in8.inv0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12870 a_22770_9598# word7.byte4.cgate0.inv1.O a_22660_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12871 VDD a_47020_4792# a_46020_4840# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12872 a_122080_3276# a_122410_3276# a_122310_3326# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X12873 a_62370_11114# word8.byte3.cgate0.inv1.O a_62260_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12874 a_65250_6462# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12875 VSS a_141060_8628# a_141020_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12876 VSS buf_in20.inv0.O buf_in20.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12877 buf_in8.inv0.O Di7 VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12878 a_49620_9714# word7.byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12879 VDD a_47020_1656# a_46020_1704# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12880 VDD buf_in1.inv0.O buf_in1.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12881 a_20820_11112# word8.byte4.tinv5.EN word8.byte4.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12882 word4.byte2.dff_7.O word4.byte2.tinv7.I VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12883 VDD buf_in23.inv0.O buf_in23.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12884 a_65250_3326# buf_in17.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12885 VSS word4.byte1.nand.B a_78780_5796# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12886 VSS word1.byte1.cgate0.nand0.B word1.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12887 VSS word7.byte1.buf_RE0.I word7.byte1.buf_RE1.I VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12888 a_166260_680# a_166050_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12889 dec8.and4_6.nand0.A A0 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12890 a_108520_6462# a_106680_6578# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12891 word1.byte4.dff_4.O word1.byte4.tinv4.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12892 a_115110_4842# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12893 a_162340_9598# a_160500_9714# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12894 word1.byte2.buf_RE1.I word1.byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12895 VSS a_62580_10088# a_62540_9598# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12896 VDD a_119640_6952# a_119600_7362# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12897 a_8370_190# word1.byte4.cgate0.inv1.O a_8260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12898 word8.byte4.tinv7.O buf_out31.inv0.I a_6420_11112# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12899 a_115830_7978# word6.byte2.dff_7.CLK a_115720_9048# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12900 word7.byte2.tinv7.O word7.byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12901 VSS a_25420_4792# a_24420_4840# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12902 a_115110_1706# buf_in12.inv1.O VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X12903 a_108520_3326# a_106680_3442# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12904 a_104640_4842# a_104410_5632# a_104080_4792# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12905 word6.byte1.tinv7.O buf_out2.inv0.I a_164100_7976# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12906 VDD word1.byte3.tinv4.I a_56820_306# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12907 a_153300_6578# word5.byte1.tinv3.EN word5.byte1.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12908 VSS word8.buf_ck1.I word8.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12909 VDD word6.byte2.tinv2.I a_110280_7976# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12910 VSS a_6420_4840# a_7980_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12911 VDD a_119640_3816# a_119600_4226# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12912 word5.byte4.tinv7.O buf_out27.inv0.I a_20820_6578# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12913 word1.byte4.tinv7.O word1.byte4.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12914 a_104640_1706# a_104410_2496# a_104080_1656# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12915 a_144340_1090# a_142500_306# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12916 word4.byte4.buf_RE0.O word4.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12917 a_11860_11114# a_10020_11112# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12918 VDD word6.byte3.cgate0.inv1.I word6.byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12919 VDD a_44580_680# a_44540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12920 VDD a_112440_8628# a_112400_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12921 VDD buf_out14.inv0.I buf_out14.inv0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X12922 word3.byte4.tinv7.O buf_out27.inv0.I a_20820_3442# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12923 VDD a_111280_7928# a_110280_7976# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12924 a_40660_5912# a_39720_4842# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12925 a_156900_7976# word6.byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12926 word2.byte4.buf_RE0.O word2.byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12927 VSS buf_out5.inv0.I buf_out5.inv0.O VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X12928 VSS buf_in25.inv0.O buf_in25.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12929 word5.byte2.dff_6.O word5.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12930 word6.byte2.tinv7.O word6.byte2.tinv3.EN a_113880_7976# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12931 VDD buf_out20.inv0.O Do19_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12932 VDD buf_in7.inv0.O buf_in7.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12933 a_159020_11114# word8.byte1.dff_7.CLK a_158850_11114# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12934 VSS a_141060_5492# word4.byte1.tinv0.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12935 VSS a_8580_11764# word8.byte4.tinv2.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12936 a_58660_9048# a_56820_7976# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12937 a_40980_5492# a_40770_4842# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12938 a_151030_6412# word5.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12939 VDD word7.byte3.tinv3.I a_53220_9714# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12940 a_11860_190# a_10020_306# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12941 word3.byte2.dff_6.O word3.byte2.tinv6.I VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12942 buf_in19.inv1.O buf_in19.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12943 a_43980_10498# a_43750_9548# a_43420_9548# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12944 word2.byte3.tinv7.O word2.byte3.buf_RE0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12945 a_119040_1090# a_118810_140# a_118480_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12946 a_44540_7362# word5.byte3.cgate0.inv1.O a_44370_6462# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12947 dec8.and4_6.nand1.OUT A2 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12948 VSS a_159060_8628# word6.byte1.tinv5.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12949 a_151030_3276# word3.byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12950 a_33420_8932# word6.byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12951 a_147330_12184# buf_in6.inv1.O VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X12952 a_58980_8628# a_58770_7978# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12953 VSS word4.buf_ck1.I word4.byte1.cgate0.nand0.B VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12954 a_19170_11114# word8.byte4.cgate0.inv1.O a_19060_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12955 a_165660_11114# a_165430_11904# a_165100_11064# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12956 a_25420_9548# word7.byte4.cgate0.inv1.O a_25650_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12957 a_123200_2776# a_122410_2496# a_123030_1706# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12958 buf_sel2.inv1.O buf_sel2.inv0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12959 word8.byte4.nand.OUT word8.byte1.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12960 a_141060_10088# a_140850_9598# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12961 a_44540_4226# word3.byte3.cgate0.inv1.O a_44370_3326# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12962 a_40150_9548# word7.byte3.cgate0.inv1.O VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X12963 word1.byte1.tinv7.O word1.byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12964 a_142500_4840# buf_out8.inv0.I word4.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12965 a_64020_3442# word3.byte3.tinv6.EN word3.byte3.tinv7.O VSS nfet_03v3 ad=357.5f pd=1.93u as=255f ps=1.45u w=850n l=300n
X12966 VSS a_12180_8628# word6.byte4.tinv3.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12967 a_101600_10498# word7.byte2.dff_7.CLK a_101430_9598# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12968 a_25420_7928# word6.byte4.cgate0.inv1.O a_25650_7978# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12969 VDD word1.buf_sel0.O word1.byte1.nand.B VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12970 a_92280_4840# word4.byte2.cgate0.latch0.I0.ENB word4.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12971 a_12180_11764# a_11970_11114# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X12972 a_147100_11064# word8.byte1.dff_7.CLK a_147330_11114# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X12973 a_126800_6462# a_126010_6412# a_126630_6462# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12974 a_159020_190# a_158230_140# a_158850_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12975 VSS a_107680_6412# a_106680_6578# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12976 a_142500_1704# buf_out8.inv0.I word2.byte1.tinv7.O VDD pfet_03v3 ad=427.5f pd=2.21u as=510f ps=2.3u w=1.7u l=300n
X12977 a_17220_9714# word7.byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12978 VSS a_44580_6952# word5.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12979 VSS word5.byte3.tinv6.I a_64020_6578# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12980 VDD a_25420_9548# a_24420_9714# VDD pfet_03v3 ad=467.5f pd=2.25u as=285f ps=1.47u w=1.705u l=300n
X12981 a_92280_1704# word2.byte2.cgate0.latch0.I0.ENB word2.byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12982 VSS a_103080_4840# a_104640_5912# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12983 VSS word8.byte1.buf_RE1.I word8.byte1.tinv7.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12984 a_126800_3326# a_126010_3276# a_126630_3326# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X12985 a_122920_4842# a_121080_4840# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12986 VDD buf_out13.inv0.O buf_out13.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X12987 VSS a_107680_3276# a_106680_3442# VSS nfet_03v3 ad=233.75f pd=1.4u as=238.325f ps=1.285u w=1000n l=300n
X12988 word6.byte4.cgate0.inv1.O word6.byte4.cgate0.inv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X12989 a_22150_140# word1.byte4.cgate0.inv1.O VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12990 word1.byte2.tinv7.O word1.byte2.tinv2.EN a_110280_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X12991 VSS a_44580_3816# word3.byte3.tinv1.I VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X12992 VDD a_55380_10088# a_55340_10498# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X12993 VSS buf_re.inv0.O buf_re.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X12994 word7.byte1.cgate0.nand0.A word7.byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X12995 VSS buf_in23.inv0.O buf_in23.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12996 VSS buf_out4.inv0.O Do3_buf VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X12997 a_122920_1706# a_121080_1704# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X12998 VSS a_146100_11112# a_147660_12184# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X12999 VDD buf_out27.inv0.O Do26_buf VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X13000 buf_in4.inv0.O Di3 VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X13001 VSS word8.byte4.inv_and.O a_36120_12068# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X13002 VSS word8.byte1.cgate0.nand0.B word8.byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X13003 a_162620_1090# word1.byte1.dff_7.CLK a_162450_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
.ends

