magic
tech gf180mcuC
timestamp 1683996514
<< nwell >>
rect 0 -9 18 57
<< properties >>
string FIXED_BBOX 0 0 18 78
<< end >>
