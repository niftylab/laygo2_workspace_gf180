magic
tech gf180mcuC
magscale 1 10
timestamp 1683398700
<< nwell >>
rect -150 -90 510 570
<< pmos >>
rect 60 136 120 476
rect 240 136 300 476
<< pdiff >>
rect -60 450 60 476
rect -60 390 -31 450
rect 31 390 60 450
rect -60 330 60 390
rect -60 270 -31 330
rect 31 270 60 330
rect -60 210 60 270
rect -60 150 -31 210
rect 31 150 60 210
rect -60 136 60 150
rect 120 450 240 476
rect 120 390 149 450
rect 211 390 240 450
rect 120 330 240 390
rect 120 270 149 330
rect 211 270 240 330
rect 120 210 240 270
rect 120 150 149 210
rect 211 150 240 210
rect 120 136 240 150
rect 300 450 420 476
rect 300 390 329 450
rect 391 390 420 450
rect 300 330 420 390
rect 300 270 329 330
rect 391 270 420 330
rect 300 210 420 270
rect 300 150 329 210
rect 391 150 420 210
rect 300 136 420 150
<< pdiffc >>
rect -31 390 31 450
rect -31 270 31 330
rect -31 150 31 210
rect 149 390 211 450
rect 149 270 211 330
rect 149 150 211 210
rect 329 390 391 450
rect 329 270 391 330
rect 329 150 391 210
<< polysilicon >>
rect 60 650 300 666
rect 60 580 150 650
rect 210 580 300 650
rect 60 566 300 580
rect 60 476 120 566
rect 240 476 300 566
rect 60 84 120 136
rect 240 84 300 136
<< polycontact >>
rect 150 580 210 650
<< metal1 >>
rect 136 650 224 672
rect 136 580 150 650
rect 210 580 224 650
rect 136 560 224 580
rect -44 450 44 476
rect -44 390 -31 450
rect 31 390 44 450
rect -44 330 44 390
rect -44 270 -31 330
rect 31 270 44 330
rect -44 210 44 270
rect -44 150 -31 210
rect 31 150 44 210
rect -44 136 44 150
rect 136 450 224 476
rect 136 390 149 450
rect 211 390 224 450
rect 136 330 224 390
rect 136 270 149 330
rect 211 270 224 330
rect 136 210 224 270
rect 136 150 149 210
rect 211 150 224 210
rect 136 136 224 150
rect 316 450 404 476
rect 316 390 329 450
rect 391 390 404 450
rect 316 330 404 390
rect 316 270 329 330
rect 391 270 404 330
rect 316 210 404 270
rect 316 150 329 210
rect 391 150 404 210
rect 316 136 404 150
<< end >>
