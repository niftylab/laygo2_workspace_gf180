magic
tech gf180mcuC
magscale 1 10
timestamp 1684460819
<< nmos >>
rect 60 306 120 476
<< ndiff >>
rect -60 459 60 476
rect -60 413 -30 459
rect 30 413 60 459
rect -60 365 60 413
rect -60 319 -30 365
rect 30 319 60 365
rect -60 306 60 319
rect 120 459 240 476
rect 120 413 150 459
rect 210 413 240 459
rect 120 365 240 413
rect 120 319 150 365
rect 210 319 240 365
rect 120 306 240 319
<< ndiffc >>
rect -30 413 30 459
rect -30 319 30 365
rect 150 413 210 459
rect 150 319 210 365
<< polysilicon >>
rect 60 650 176 666
rect 60 580 110 650
rect 160 580 176 650
rect 60 566 176 580
rect 60 476 120 566
rect 60 262 120 306
<< polycontact >>
rect 110 580 160 650
<< metal1 >>
rect 94 650 224 672
rect 94 580 110 650
rect 160 580 224 650
rect 94 560 224 580
rect -44 459 44 476
rect -44 413 -30 459
rect 30 413 44 459
rect -44 365 44 413
rect -44 319 -30 365
rect 30 319 44 365
rect -44 280 44 319
rect 136 459 224 476
rect 136 413 150 459
rect 210 413 224 459
rect 136 365 224 413
rect 136 319 150 365
rect 210 319 224 365
rect 136 280 224 319
<< end >>
