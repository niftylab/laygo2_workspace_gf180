magic
tech gf180mcuC
magscale 1 10
timestamp 1689441100
<< nwell >>
rect 0 990 2700 1660
<< nmos >>
rect 220 190 280 360
rect 390 190 450 360
rect 550 190 610 360
rect 720 190 780 360
rect 830 190 890 360
rect 1000 190 1060 360
rect 1110 190 1170 360
rect 1280 190 1340 360
rect 1390 190 1450 360
rect 1560 190 1620 360
rect 1880 190 1940 360
rect 2200 190 2260 360
rect 2370 190 2430 360
<< pmos >>
rect 220 1090 280 1430
rect 390 1090 450 1430
rect 550 1090 610 1430
rect 720 1090 780 1430
rect 830 1090 890 1430
rect 1000 1090 1060 1430
rect 1110 1090 1170 1430
rect 1280 1090 1340 1430
rect 1390 1090 1450 1430
rect 1560 1090 1620 1430
rect 1880 1090 1940 1430
rect 2200 1090 2260 1430
rect 2370 1090 2430 1430
<< ndiff >>
rect 120 298 220 360
rect 120 252 142 298
rect 188 252 220 298
rect 120 190 220 252
rect 280 298 390 360
rect 280 252 312 298
rect 358 252 390 298
rect 280 190 390 252
rect 450 190 550 360
rect 610 298 720 360
rect 610 252 642 298
rect 688 252 720 298
rect 610 190 720 252
rect 780 190 830 360
rect 890 258 1000 360
rect 890 212 922 258
rect 968 212 1000 258
rect 890 190 1000 212
rect 1060 190 1110 360
rect 1170 298 1280 360
rect 1170 252 1202 298
rect 1248 252 1280 298
rect 1170 190 1280 252
rect 1340 190 1390 360
rect 1450 298 1560 360
rect 1450 252 1482 298
rect 1528 252 1560 298
rect 1450 190 1560 252
rect 1620 298 1720 360
rect 1620 252 1652 298
rect 1698 252 1720 298
rect 1620 190 1720 252
rect 1780 263 1880 360
rect 1780 217 1802 263
rect 1848 217 1880 263
rect 1780 190 1880 217
rect 1940 298 2040 360
rect 1940 252 1972 298
rect 2018 252 2040 298
rect 1940 190 2040 252
rect 2100 298 2200 360
rect 2100 252 2122 298
rect 2168 252 2200 298
rect 2100 190 2200 252
rect 2260 298 2370 360
rect 2260 252 2292 298
rect 2338 252 2370 298
rect 2260 190 2370 252
rect 2430 298 2530 360
rect 2430 252 2462 298
rect 2508 252 2530 298
rect 2430 190 2530 252
<< pdiff >>
rect 120 1377 220 1430
rect 120 1143 142 1377
rect 188 1143 220 1377
rect 120 1090 220 1143
rect 280 1377 390 1430
rect 280 1143 312 1377
rect 358 1143 390 1377
rect 280 1090 390 1143
rect 450 1090 550 1430
rect 610 1377 720 1430
rect 610 1143 642 1377
rect 688 1143 720 1377
rect 610 1090 720 1143
rect 780 1090 830 1430
rect 890 1377 1000 1430
rect 890 1143 922 1377
rect 968 1143 1000 1377
rect 890 1090 1000 1143
rect 1060 1090 1110 1430
rect 1170 1405 1280 1430
rect 1170 1265 1202 1405
rect 1248 1265 1280 1405
rect 1170 1090 1280 1265
rect 1340 1090 1390 1430
rect 1450 1405 1560 1430
rect 1450 1265 1482 1405
rect 1528 1265 1560 1405
rect 1450 1090 1560 1265
rect 1620 1377 1720 1430
rect 1620 1143 1652 1377
rect 1698 1143 1720 1377
rect 1620 1090 1720 1143
rect 1780 1377 1880 1430
rect 1780 1143 1802 1377
rect 1848 1143 1880 1377
rect 1780 1090 1880 1143
rect 1940 1377 2040 1430
rect 1940 1143 1972 1377
rect 2018 1143 2040 1377
rect 1940 1090 2040 1143
rect 2100 1377 2200 1430
rect 2100 1143 2122 1377
rect 2168 1143 2200 1377
rect 2100 1090 2200 1143
rect 2260 1377 2370 1430
rect 2260 1143 2292 1377
rect 2338 1143 2370 1377
rect 2260 1090 2370 1143
rect 2430 1377 2530 1430
rect 2430 1143 2462 1377
rect 2508 1143 2530 1377
rect 2430 1090 2530 1143
<< ndiffc >>
rect 142 252 188 298
rect 312 252 358 298
rect 642 252 688 298
rect 922 212 968 258
rect 1202 252 1248 298
rect 1482 252 1528 298
rect 1652 252 1698 298
rect 1802 217 1848 263
rect 1972 252 2018 298
rect 2122 252 2168 298
rect 2292 252 2338 298
rect 2462 252 2508 298
<< pdiffc >>
rect 142 1143 188 1377
rect 312 1143 358 1377
rect 642 1143 688 1377
rect 922 1143 968 1377
rect 1202 1265 1248 1405
rect 1482 1265 1528 1405
rect 1652 1143 1698 1377
rect 1802 1143 1848 1377
rect 1972 1143 2018 1377
rect 2122 1143 2168 1377
rect 2292 1143 2338 1377
rect 2462 1143 2508 1377
<< psubdiff >>
rect 120 98 210 120
rect 120 52 142 98
rect 188 52 210 98
rect 120 30 210 52
rect 360 98 450 120
rect 360 52 382 98
rect 428 52 450 98
rect 360 30 450 52
rect 600 98 690 120
rect 600 52 622 98
rect 668 52 690 98
rect 600 30 690 52
rect 840 98 930 120
rect 840 52 862 98
rect 908 52 930 98
rect 840 30 930 52
rect 1080 98 1170 120
rect 1080 52 1102 98
rect 1148 52 1170 98
rect 1080 30 1170 52
rect 1320 98 1410 120
rect 1320 52 1342 98
rect 1388 52 1410 98
rect 1320 30 1410 52
rect 1560 98 1650 120
rect 1560 52 1582 98
rect 1628 52 1650 98
rect 1560 30 1650 52
rect 1800 98 1890 120
rect 1800 52 1822 98
rect 1868 52 1890 98
rect 1800 30 1890 52
rect 2040 98 2130 120
rect 2040 52 2062 98
rect 2108 52 2130 98
rect 2040 30 2130 52
rect 2280 98 2370 120
rect 2280 52 2302 98
rect 2348 52 2370 98
rect 2280 30 2370 52
<< nsubdiff >>
rect 120 1568 210 1590
rect 120 1522 142 1568
rect 188 1522 210 1568
rect 120 1500 210 1522
rect 360 1568 450 1590
rect 360 1522 382 1568
rect 428 1522 450 1568
rect 360 1500 450 1522
rect 600 1568 690 1590
rect 600 1522 622 1568
rect 668 1522 690 1568
rect 600 1500 690 1522
rect 840 1568 930 1590
rect 840 1522 862 1568
rect 908 1522 930 1568
rect 840 1500 930 1522
rect 1080 1568 1170 1590
rect 1080 1522 1102 1568
rect 1148 1522 1170 1568
rect 1080 1500 1170 1522
rect 1320 1568 1410 1590
rect 1320 1522 1342 1568
rect 1388 1522 1410 1568
rect 1320 1500 1410 1522
rect 1560 1568 1650 1590
rect 1560 1522 1582 1568
rect 1628 1522 1650 1568
rect 1560 1500 1650 1522
rect 1800 1568 1890 1590
rect 1800 1522 1822 1568
rect 1868 1522 1890 1568
rect 1800 1500 1890 1522
rect 2040 1568 2130 1590
rect 2040 1522 2062 1568
rect 2108 1522 2130 1568
rect 2040 1500 2130 1522
rect 2280 1568 2370 1590
rect 2280 1522 2302 1568
rect 2348 1522 2370 1568
rect 2280 1500 2370 1522
<< psubdiffcont >>
rect 142 52 188 98
rect 382 52 428 98
rect 622 52 668 98
rect 862 52 908 98
rect 1102 52 1148 98
rect 1342 52 1388 98
rect 1582 52 1628 98
rect 1822 52 1868 98
rect 2062 52 2108 98
rect 2302 52 2348 98
<< nsubdiffcont >>
rect 142 1522 188 1568
rect 382 1522 428 1568
rect 622 1522 668 1568
rect 862 1522 908 1568
rect 1102 1522 1148 1568
rect 1342 1522 1388 1568
rect 1582 1522 1628 1568
rect 1822 1522 1868 1568
rect 2062 1522 2108 1568
rect 2302 1522 2348 1568
<< polysilicon >>
rect 220 1430 280 1480
rect 390 1430 450 1480
rect 550 1430 610 1480
rect 720 1430 780 1480
rect 830 1430 890 1480
rect 1000 1430 1060 1480
rect 1110 1430 1170 1480
rect 1280 1430 1340 1480
rect 1390 1430 1450 1480
rect 1560 1430 1620 1480
rect 1880 1430 1940 1480
rect 2200 1430 2260 1480
rect 2370 1430 2430 1480
rect 220 910 280 1090
rect 220 883 340 910
rect 220 837 267 883
rect 313 837 340 883
rect 220 810 340 837
rect 220 360 280 810
rect 390 780 450 1090
rect 550 910 610 1090
rect 550 883 650 910
rect 550 837 577 883
rect 623 837 650 883
rect 550 810 650 837
rect 390 753 510 780
rect 390 707 437 753
rect 483 707 510 753
rect 390 680 510 707
rect 390 360 450 680
rect 720 640 780 1090
rect 830 1040 890 1090
rect 1000 1040 1060 1090
rect 830 1013 1060 1040
rect 830 970 867 1013
rect 840 967 867 970
rect 913 970 1060 1013
rect 913 967 940 970
rect 840 920 940 967
rect 1110 640 1170 1090
rect 1280 910 1340 1090
rect 1240 883 1340 910
rect 1240 837 1267 883
rect 1313 837 1340 883
rect 1240 810 1340 837
rect 1390 780 1450 1090
rect 1560 910 1620 1090
rect 1560 883 1660 910
rect 1560 837 1587 883
rect 1633 837 1660 883
rect 1560 810 1660 837
rect 1380 753 1490 780
rect 1380 707 1407 753
rect 1453 707 1490 753
rect 1380 680 1490 707
rect 1240 640 1340 650
rect 550 623 1340 640
rect 550 580 1267 623
rect 550 360 610 580
rect 1240 577 1267 580
rect 1313 577 1340 623
rect 1240 550 1340 577
rect 680 493 780 520
rect 840 500 940 520
rect 680 447 707 493
rect 753 447 780 493
rect 680 420 780 447
rect 720 360 780 420
rect 830 493 1060 500
rect 830 447 867 493
rect 913 447 1060 493
rect 830 420 1060 447
rect 830 360 890 420
rect 1000 360 1060 420
rect 1110 483 1210 510
rect 1110 437 1137 483
rect 1183 437 1210 483
rect 1110 410 1210 437
rect 1110 360 1170 410
rect 1280 360 1340 550
rect 1390 360 1450 680
rect 1560 360 1620 810
rect 1880 650 1940 1090
rect 2200 650 2260 1090
rect 2370 910 2430 1090
rect 2310 883 2430 910
rect 2310 837 2337 883
rect 2383 837 2430 883
rect 2310 810 2430 837
rect 1820 623 1940 650
rect 1820 577 1847 623
rect 1893 577 1940 623
rect 1820 550 1940 577
rect 2140 623 2260 650
rect 2140 577 2187 623
rect 2233 577 2260 623
rect 2140 550 2260 577
rect 1880 360 1940 550
rect 2200 360 2260 550
rect 2370 360 2430 810
rect 220 140 280 190
rect 390 140 450 190
rect 550 140 610 190
rect 720 140 780 190
rect 830 140 890 190
rect 1000 140 1060 190
rect 1110 140 1170 190
rect 1280 140 1340 190
rect 1390 140 1450 190
rect 1560 140 1620 190
rect 1880 140 1940 190
rect 2200 140 2260 190
rect 2370 140 2430 190
<< polycontact >>
rect 267 837 313 883
rect 577 837 623 883
rect 437 707 483 753
rect 867 967 913 1013
rect 1267 837 1313 883
rect 1587 837 1633 883
rect 1407 707 1453 753
rect 1267 577 1313 623
rect 707 447 753 493
rect 867 447 913 493
rect 1137 437 1183 483
rect 2337 837 2383 883
rect 1847 577 1893 623
rect 2187 577 2233 623
<< metal1 >>
rect 110 1610 2540 1630
rect 110 1568 280 1610
rect 390 1568 580 1610
rect 690 1568 880 1610
rect 990 1568 1180 1610
rect 110 1522 142 1568
rect 188 1522 280 1568
rect 428 1522 580 1568
rect 690 1522 862 1568
rect 990 1522 1102 1568
rect 1148 1522 1180 1568
rect 110 1520 280 1522
rect 390 1520 580 1522
rect 690 1520 880 1522
rect 990 1520 1180 1522
rect 1290 1568 1480 1610
rect 1590 1568 1780 1610
rect 1890 1568 2080 1610
rect 1290 1522 1342 1568
rect 1388 1522 1480 1568
rect 1628 1522 1780 1568
rect 1890 1522 2062 1568
rect 1290 1520 1480 1522
rect 1590 1520 1780 1522
rect 1890 1520 2080 1522
rect 2190 1520 2290 1610
rect 2400 1520 2540 1610
rect 110 1500 2540 1520
rect 140 1377 190 1430
rect 140 1143 142 1377
rect 188 1143 190 1377
rect 140 520 190 1143
rect 310 1377 360 1500
rect 310 1143 312 1377
rect 358 1143 360 1377
rect 310 1090 360 1143
rect 640 1377 690 1430
rect 640 1143 642 1377
rect 688 1143 690 1377
rect 640 1040 690 1143
rect 920 1377 970 1500
rect 920 1143 922 1377
rect 968 1143 970 1377
rect 1200 1405 1250 1430
rect 1200 1265 1202 1405
rect 1248 1265 1250 1405
rect 1200 1240 1250 1265
rect 1480 1405 1530 1500
rect 1480 1265 1482 1405
rect 1528 1265 1530 1405
rect 1480 1240 1530 1265
rect 1650 1377 1700 1430
rect 920 1090 970 1143
rect 1020 1190 1250 1240
rect 310 990 690 1040
rect 840 1013 940 1020
rect 310 890 360 990
rect 840 967 867 1013
rect 913 967 940 1013
rect 840 960 940 967
rect 240 883 360 890
rect 240 837 267 883
rect 313 837 360 883
rect 240 830 360 837
rect 550 886 780 890
rect 550 883 704 886
rect 550 837 577 883
rect 623 837 704 883
rect 550 834 704 837
rect 756 834 780 886
rect 550 830 780 834
rect 130 496 190 520
rect 130 444 134 496
rect 186 444 190 496
rect 310 500 360 830
rect 410 756 510 760
rect 410 704 434 756
rect 486 704 510 756
rect 410 700 510 704
rect 700 500 760 830
rect 860 500 920 960
rect 1020 740 1070 1190
rect 1650 1143 1652 1377
rect 1698 1143 1700 1377
rect 1370 1016 1470 1020
rect 1370 964 1394 1016
rect 1446 964 1470 1016
rect 1370 960 1470 964
rect 1650 1000 1700 1143
rect 1800 1377 1850 1500
rect 1800 1143 1802 1377
rect 1848 1143 1850 1377
rect 1800 1090 1850 1143
rect 1970 1377 2020 1430
rect 1970 1143 1972 1377
rect 2018 1143 2020 1377
rect 1010 690 1070 740
rect 1130 886 1340 890
rect 1130 834 1264 886
rect 1316 834 1340 886
rect 1130 830 1340 834
rect 310 450 510 500
rect 130 420 190 444
rect 140 298 190 420
rect 430 360 510 450
rect 680 493 780 500
rect 680 447 707 493
rect 753 447 780 493
rect 680 440 780 447
rect 840 496 940 500
rect 840 444 864 496
rect 916 444 940 496
rect 840 440 940 444
rect 1010 370 1060 690
rect 1130 490 1190 830
rect 1390 760 1450 960
rect 1650 950 1810 1000
rect 1560 886 1660 890
rect 1560 834 1584 886
rect 1636 834 1660 886
rect 1560 830 1660 834
rect 1750 760 1810 950
rect 1380 756 1490 760
rect 1380 704 1404 756
rect 1456 704 1490 756
rect 1380 700 1490 704
rect 1650 710 1810 760
rect 1390 690 1470 700
rect 1240 626 1340 630
rect 1240 574 1264 626
rect 1316 574 1340 626
rect 1240 570 1340 574
rect 1650 626 1710 710
rect 1840 630 1900 650
rect 1970 630 2020 1143
rect 2120 1377 2170 1430
rect 2120 1143 2122 1377
rect 2168 1143 2170 1377
rect 2120 890 2170 1143
rect 2290 1377 2340 1500
rect 2290 1143 2292 1377
rect 2338 1143 2340 1377
rect 2290 1090 2340 1143
rect 2460 1377 2510 1430
rect 2460 1143 2462 1377
rect 2508 1143 2510 1377
rect 2460 1030 2510 1143
rect 2460 1016 2560 1030
rect 2460 964 2484 1016
rect 2536 964 2560 1016
rect 2460 960 2560 964
rect 2460 950 2550 960
rect 2120 883 2410 890
rect 2120 837 2337 883
rect 2383 837 2410 883
rect 2120 830 2410 837
rect 1650 574 1654 626
rect 1706 574 1710 626
rect 1650 550 1710 574
rect 1820 623 1920 630
rect 1820 577 1847 623
rect 1893 577 1920 623
rect 1820 570 1920 577
rect 1970 626 2260 630
rect 1970 574 2184 626
rect 2236 574 2260 626
rect 1970 570 2260 574
rect 1110 483 1210 490
rect 1110 437 1137 483
rect 1183 437 1210 483
rect 1110 430 1210 437
rect 1010 366 1280 370
rect 140 252 142 298
rect 188 252 190 298
rect 140 190 190 252
rect 310 298 360 360
rect 430 310 690 360
rect 1010 320 1204 366
rect 310 252 312 298
rect 358 252 360 298
rect 310 120 360 252
rect 640 298 690 310
rect 640 252 642 298
rect 688 252 690 298
rect 1200 314 1204 320
rect 1256 314 1280 366
rect 1200 310 1280 314
rect 1200 298 1250 310
rect 640 190 690 252
rect 920 258 970 280
rect 920 212 922 258
rect 968 212 970 258
rect 920 120 970 212
rect 1200 252 1202 298
rect 1248 252 1250 298
rect 1200 190 1250 252
rect 1480 298 1530 360
rect 1480 252 1482 298
rect 1528 252 1530 298
rect 1480 120 1530 252
rect 1650 298 1700 550
rect 1840 400 1900 570
rect 1820 396 1920 400
rect 1820 344 1844 396
rect 1896 344 1920 396
rect 1820 340 1920 344
rect 1650 252 1652 298
rect 1698 252 1700 298
rect 1970 298 2020 570
rect 2340 500 2390 830
rect 2290 477 2390 500
rect 2290 460 2310 477
rect 1650 190 1700 252
rect 1800 263 1850 290
rect 1800 217 1802 263
rect 1848 217 1850 263
rect 1800 120 1850 217
rect 1970 252 1972 298
rect 2018 252 2020 298
rect 1970 190 2020 252
rect 2120 425 2310 460
rect 2370 425 2390 477
rect 2120 410 2390 425
rect 2120 298 2170 410
rect 2120 252 2122 298
rect 2168 252 2170 298
rect 2120 190 2170 252
rect 2290 298 2340 360
rect 2290 252 2292 298
rect 2338 252 2340 298
rect 2290 120 2340 252
rect 2460 298 2510 950
rect 2460 252 2462 298
rect 2508 252 2510 298
rect 2460 190 2510 252
rect 110 98 2520 120
rect 110 52 142 98
rect 188 60 382 98
rect 428 60 622 98
rect 668 60 862 98
rect 908 60 1102 98
rect 1148 60 1342 98
rect 1388 60 1582 98
rect 1628 60 1822 98
rect 1868 60 2062 98
rect 2108 60 2302 98
rect 2348 60 2520 98
rect 188 52 310 60
rect 428 52 530 60
rect 668 52 780 60
rect 908 52 1030 60
rect 1148 52 1280 60
rect 110 -30 310 52
rect 420 -30 530 52
rect 640 -30 780 52
rect 890 -30 1030 52
rect 1140 -30 1280 52
rect 1390 -30 1530 60
rect 1640 -30 1780 60
rect 1890 -30 2030 60
rect 2140 -30 2280 60
rect 2390 -30 2520 60
rect 110 -60 2520 -30
<< via1 >>
rect 280 1568 390 1610
rect 580 1568 690 1610
rect 880 1568 990 1610
rect 280 1522 382 1568
rect 382 1522 390 1568
rect 580 1522 622 1568
rect 622 1522 668 1568
rect 668 1522 690 1568
rect 880 1522 908 1568
rect 908 1522 990 1568
rect 280 1520 390 1522
rect 580 1520 690 1522
rect 880 1520 990 1522
rect 1180 1520 1290 1610
rect 1480 1568 1590 1610
rect 1780 1568 1890 1610
rect 2080 1568 2190 1610
rect 1480 1522 1582 1568
rect 1582 1522 1590 1568
rect 1780 1522 1822 1568
rect 1822 1522 1868 1568
rect 1868 1522 1890 1568
rect 2080 1522 2108 1568
rect 2108 1522 2190 1568
rect 1480 1520 1590 1522
rect 1780 1520 1890 1522
rect 2080 1520 2190 1522
rect 2290 1568 2400 1610
rect 2290 1522 2302 1568
rect 2302 1522 2348 1568
rect 2348 1522 2400 1568
rect 2290 1520 2400 1522
rect 704 834 756 886
rect 134 444 186 496
rect 434 753 486 756
rect 434 707 437 753
rect 437 707 483 753
rect 483 707 486 753
rect 434 704 486 707
rect 1394 964 1446 1016
rect 1264 883 1316 886
rect 1264 837 1267 883
rect 1267 837 1313 883
rect 1313 837 1316 883
rect 1264 834 1316 837
rect 864 493 916 496
rect 864 447 867 493
rect 867 447 913 493
rect 913 447 916 493
rect 864 444 916 447
rect 1584 883 1636 886
rect 1584 837 1587 883
rect 1587 837 1633 883
rect 1633 837 1636 883
rect 1584 834 1636 837
rect 1404 753 1456 756
rect 1404 707 1407 753
rect 1407 707 1453 753
rect 1453 707 1456 753
rect 1404 704 1456 707
rect 1264 623 1316 626
rect 1264 577 1267 623
rect 1267 577 1313 623
rect 1313 577 1316 623
rect 1264 574 1316 577
rect 2484 964 2536 1016
rect 1654 574 1706 626
rect 2184 623 2236 626
rect 2184 577 2187 623
rect 2187 577 2233 623
rect 2233 577 2236 623
rect 2184 574 2236 577
rect 1204 314 1256 366
rect 1844 344 1896 396
rect 2310 425 2370 477
rect 310 52 382 60
rect 382 52 420 60
rect 530 52 622 60
rect 622 52 640 60
rect 780 52 862 60
rect 862 52 890 60
rect 1030 52 1102 60
rect 1102 52 1140 60
rect 1280 52 1342 60
rect 1342 52 1388 60
rect 1388 52 1390 60
rect 310 -30 420 52
rect 530 -30 640 52
rect 780 -30 890 52
rect 1030 -30 1140 52
rect 1280 -30 1390 52
rect 1530 52 1582 60
rect 1582 52 1628 60
rect 1628 52 1640 60
rect 1530 -30 1640 52
rect 1780 52 1822 60
rect 1822 52 1868 60
rect 1868 52 1890 60
rect 1780 -30 1890 52
rect 2030 52 2062 60
rect 2062 52 2108 60
rect 2108 52 2140 60
rect 2030 -30 2140 52
rect 2280 52 2302 60
rect 2302 52 2348 60
rect 2348 52 2390 60
rect 2280 -30 2390 52
<< metal2 >>
rect 0 1610 2650 1654
rect 0 1520 280 1610
rect 390 1520 580 1610
rect 690 1520 880 1610
rect 990 1520 1180 1610
rect 1290 1520 1480 1610
rect 1590 1520 1780 1610
rect 1890 1520 2080 1610
rect 2190 1520 2290 1610
rect 2400 1520 2650 1610
rect 0 1480 2650 1520
rect 1380 1020 1460 1030
rect 2470 1020 2550 1030
rect 1370 1016 2010 1020
rect 1370 964 1394 1016
rect 1446 964 2010 1016
rect 1370 960 2010 964
rect 2110 960 2120 1020
rect 2200 1016 2560 1020
rect 2200 964 2484 1016
rect 2536 964 2560 1016
rect 2200 960 2560 964
rect 1380 950 1460 960
rect 680 890 770 900
rect 1240 890 1340 900
rect 1570 890 1650 900
rect 760 886 1660 890
rect 760 834 1264 886
rect 1316 834 1584 886
rect 1636 834 1660 886
rect 760 830 1660 834
rect 680 820 770 830
rect 1240 820 1340 830
rect 1570 820 1650 830
rect 320 690 330 770
rect 400 760 510 770
rect 1390 760 1470 770
rect 400 756 540 760
rect 400 704 434 756
rect 486 704 540 756
rect 400 700 540 704
rect 1380 756 1480 760
rect 1380 704 1404 756
rect 1456 704 1480 756
rect 1380 700 1480 704
rect 400 690 510 700
rect 1390 690 1470 700
rect 1250 630 1330 640
rect 1640 630 1720 640
rect 1950 630 2010 960
rect 2470 950 2550 960
rect 2170 630 2250 640
rect 1240 626 1740 630
rect 1240 574 1264 626
rect 1316 574 1654 626
rect 1706 574 1740 626
rect 1240 570 1740 574
rect 1950 626 2260 630
rect 1950 574 2184 626
rect 2236 574 2260 626
rect 1950 570 2260 574
rect 1250 560 1330 570
rect 1640 560 1720 570
rect 2170 560 2250 570
rect 120 500 200 510
rect 850 500 930 510
rect 120 496 940 500
rect 120 444 134 496
rect 186 444 864 496
rect 916 444 940 496
rect 120 440 940 444
rect 2110 479 2390 480
rect 120 430 200 440
rect 850 430 930 440
rect 2110 423 2310 479
rect 2370 423 2390 479
rect 2110 420 2390 423
rect 1830 400 1910 410
rect 1730 396 1920 400
rect 1190 370 1270 380
rect 1730 370 1844 396
rect 1180 366 1844 370
rect 1180 314 1204 366
rect 1256 344 1844 366
rect 1896 344 1920 396
rect 1256 340 1920 344
rect 1256 330 1910 340
rect 1256 314 1790 330
rect 1180 310 1790 314
rect 1190 300 1270 310
rect 0 60 2680 90
rect 0 -30 310 60
rect 420 -30 530 60
rect 640 -30 780 60
rect 890 -30 1030 60
rect 1140 -30 1280 60
rect 1390 -30 1530 60
rect 1640 -30 1780 60
rect 1890 -30 2030 60
rect 2140 -30 2280 60
rect 2390 -30 2680 60
rect 0 -80 2680 -30
<< via2 >>
rect 2120 960 2200 1020
rect 680 886 760 890
rect 680 834 704 886
rect 704 834 756 886
rect 756 834 760 886
rect 680 830 760 834
rect 330 690 400 770
rect 2310 477 2370 479
rect 2310 425 2370 477
rect 2310 423 2370 425
<< metal3 >>
rect 2116 1020 2204 1140
rect 2116 960 2120 1020
rect 2200 960 2204 1020
rect 316 770 404 952
rect 316 690 330 770
rect 400 690 404 770
rect 316 616 404 690
rect 676 890 764 952
rect 676 830 680 890
rect 760 830 764 890
rect 676 616 764 830
rect 2116 420 2204 960
rect 2290 479 2390 1140
rect 2290 423 2310 479
rect 2370 423 2390 479
rect 2290 420 2390 423
<< labels >>
rlabel metal1 2120 830 2410 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.QN
rlabel metal1 2340 410 2390 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.QN
rlabel metal1 2120 410 2390 460 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.QN
rlabel metal1 2120 830 2170 1430 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.QN
rlabel metal1 2120 190 2170 460 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.QN
rlabel metal1 2460 960 2560 1030 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel metal1 2460 950 2550 1030 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel metal1 2460 190 2510 1430 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel metal2 2460 960 2560 1020 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel metal2 2470 950 2550 1030 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel metal2 410 700 510 760 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.D
rlabel metal2 380 700 540 760 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.D
rlabel metal2 410 690 510 770 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.D
rlabel metal2 1560 830 1660 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal2 1130 830 1340 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal1 1110 430 1210 490 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal1 1130 430 1190 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal1 550 830 780 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal1 680 440 780 500 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal1 700 440 760 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel space 680 830 1660 890 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal2 1570 820 1650 900 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel metal2 1240 820 1340 900 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel space 680 820 770 900 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel via1 704 834 756 886 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel via1 1264 834 1316 886 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel space 2290 0 2340 360 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel space 1800 0 1850 290 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel metal1 1480 0 1530 360 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel metal1 920 0 970 280 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel metal1 1480 1240 1530 1620 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel metal1 920 1090 970 1620 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel metal1 310 0 360 360 4 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel metal1 310 1090 360 1620 4 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel via1 1584 834 1636 886 4 gf180mcu_osu_sc_gp12t3v3__dff_1_0.CLK
rlabel via1 2484 964 2536 1016 4 gf180mcu_osu_sc_gp12t3v3__dff_1_0.Q
rlabel via1 434 704 486 756 4 gf180mcu_osu_sc_gp12t3v3__dff_1_0.D
rlabel space 30 0 2630 120 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VSS
rlabel nwell 1800 1090 1850 1620 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel nwell 2290 1090 2340 1620 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel nwell 30 1500 2630 1620 1 gf180mcu_osu_sc_gp12t3v3__dff_1_0.VDD
rlabel metal3 316 616 400 950 1 I
port 1 n
rlabel metal3 676 616 760 950 1 CLK
port 2 n
rlabel metal3 2116 420 2200 1140 1 O
port 3 n
rlabel metal3 2290 430 2390 1140 1 O_bar
port 4 n
rlabel metal2 0 -80 2670 80 1 VSS
port 6 n
rlabel metal2 10 1520 2640 1640 1 VDD
port 5 n
<< end >>
