** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/clk_gate.sch
.subckt clk_gate CK_I VDD VSS EN CK_O
*.PININFO CK_I:I VDD:B VSS:B EN:I CK_O:O
X_inv1 CK_I VDD VSS net1 inv NF=NF
X_latch1 EN net1 CK_I VSS VDD net2 latch NF=NF
X_nand1 CK_I net2 net3 VDD VSS nand NF=NF
X_inv2 net3 VDD VSS CK_O inv NF=NF*3
.ends

* expanding   symbol:  xschem_lib/DFFRAM_full_custom/inv.sym # of pins=4
** sym_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/inv.sym
** sch_path: /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/inv.sch
.subckt inv  X VDD VSS Y   NF=2
*.PININFO VSS:B X:I Y:O VDD:B
XM1 Y X VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y X VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/latch.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/latch.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/latch.sch
.subckt latch  IN CLK CLKB VSS VDD OUT   NF=2
*.PININFO CLKB:I IN:I CLK:I VDD:B VSS:B OUT:O
X_tinv1 IN CLK CLKB VDD VSS net1 tinv NF=NF
X_inv1 net1 VDD VSS OUT inv NF=NF
X_tinv_small1 OUT CLKB CLK VDD VSS net1 tinv_small
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/nand.sym # of pins=5
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nand.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/nand.sch
.subckt nand  B A Y VDD VSS   NF=2
*.PININFO Y:O A:I VDD:B VSS:B B:I
XM2 net1 B VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y B VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 Y A VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 Y A net1 VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/tinv.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv.sch
.subckt tinv  X EN ENB VDD VSS Y   NF=2
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y ENB net2 VDD pfet_03v3 L=0.28u W=NF*1.7u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y EN net1 VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 X VSS VSS nfet_03v3 L=0.28u W=NF*0.85u nf=NF ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  xschem_lib/DFFRAM_full_custom/tinv_small.sym # of pins=6
** sym_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv_small.sym
** sch_path:
*+ /home/sonic/gf180_tutorial/laygo2_workspace_gf180/xschem_lib/DFFRAM_full_custom/tinv_small.sch
.subckt tinv_small  X EN ENB VDD VSS Y
*.PININFO X:I ENB:I EN:I Y:O VDD:B VSS:B
XM1 net2 X VDD VDD pfet_03v3 L=0.28u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 Y ENB net2 VDD pfet_03v3 L=0.28u W=1.7u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 Y EN net1 VSS nfet_03v3 L=0.28u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 net1 X VSS VSS nfet_03v3 L=0.28u W=0.85u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.end
