* NGSPICE file created from word_flat.ext - technology: gf180mcuC

.subckt word_flat SEL WE3 WE2 WE1 WE0 CLK RE Do24 Di24 Do25 Di25 Do26 Di26 Do27 Di27
+ Do28 Di28 Do29 Di29 Do30 Di30 Do31 Di31 Do16 Di16 Do17 Di17 Do18 Di18 Do19 Di19
+ Do20 Di20 Do21 Di21 Do22 Di22 Do23 Di23 Do8 Di8 Do9 Di9 Do10 Di10 Do11 Di11 Do12
+ Di12 Do13 Di13 Do14 Di14 Do15 Di15 Do0 Di0 Do1 Di1 Do2 Di2 Do3 Di3 Do4 Di4 Do5 Di5
+ Do6 Di6 Do7 Di7 VDD VSS
X0 a_15900_190# byte4.dff_4.CLK a_15340_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1 a_130770_190# byte2.dff_7.CLK a_130660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X2 a_1380_680# a_1170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X3 VDD byte4.cgate0.nand0.A a_37200_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X4 a_37560_306# byte4.cgate0.latch0.I0.O byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X5 VDD byte3.cgate0.latch0.I0.I a_78600_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X6 buf_sel1.O buf_sel1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X7 VSS a_1380_680# byte4.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X8 byte4.inv_and.O byte4.inv_and.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X9 VSS a_42420_680# byte3.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X10 a_20070_190# a_19450_140# a_19960_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X11 byte3.dff_5.O byte3.dff_5.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X12 Do14 byte2.tinv1.ENB a_109740_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X13 VSS a_159240_190# a_159900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X14 VDD byte3.buf_RE1.I byte3.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X15 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X16 byte2.dff_2.O byte2.dff_2.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X17 a_166900_140# a_167230_140# a_167130_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X18 a_171520_190# a_170580_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X19 a_64890_190# a_64270_140# a_64780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X20 a_144550_140# byte1.dff_0.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X21 a_62760_1092# byte3.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X22 VDD byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X23 VDD byte2.tinv5.I a_124860_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X24 byte4.buf_RE0.O byte4.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X25 a_46200_680# a_45990_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X26 byte2.dff_5.O byte2.dff_5.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X27 a_155890_140# byte1.dff_3.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X28 VDD a_8940_680# a_8900_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X29 a_23130_190# Di25 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X30 VSS byte2.buf_RE0.I byte2.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X31 byte4.cgate0.nand0.OUT byte4.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X32 a_152620_1090# a_151680_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X33 a_45270_1090# Di22 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X34 a_49980_680# a_49770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X35 a_4230_190# Di30 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X36 a_55200_1092# byte3.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X37 a_57330_190# a_56710_140# a_57220_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X38 VDD byte2.cgate0.latch0.I0.O byte2.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X39 byte2.inv_and.O byte2.inv_and.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X40 VSS a_110820_190# a_111480_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X41 a_154380_306# byte1.tinv2.EN Do5 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X42 a_146820_1092# byte1.tinv0.ENB Do7 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X43 byte4.inv_and.O byte4.inv_and.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X44 VSS byte4.inv_and.I byte4.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X45 a_61320_680# a_61110_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X46 VDD a_151780_140# a_151680_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X47 byte4.dff_4.O byte4.dff_4.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X48 VDD a_46200_680# byte3.dff_1.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X49 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X50 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X51 VDD a_144120_190# a_144780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X52 a_56610_190# Di19 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X53 a_107700_1090# a_107470_140# a_107140_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X54 a_27240_1090# a_27010_140# a_26680_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X55 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X56 VDD byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X57 a_17940_1092# byte4.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X58 a_152340_190# byte1.dff_2.CLK a_151780_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X59 a_53550_190# byte3.dff_3.CLK a_53440_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X60 Do15 byte2.tinv0.EN a_105960_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X61 VDD a_166800_190# a_167460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X62 a_163680_190# byte1.dff_5.CLK a_163120_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X63 a_64890_190# byte3.dff_6.CLK a_64780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X64 byte3.buf_RE0.O byte3.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X65 VSS a_118380_190# a_119040_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X66 a_19120_140# byte4.dff_5.CLK a_19350_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X67 byte4.nand.OUT byte4.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X68 a_61280_1090# byte3.dff_5.CLK a_61110_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X69 a_68880_680# a_68670_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X70 a_145060_190# a_144120_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X71 byte4.dff_6.O byte4.dff_6.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X72 VSS a_46200_680# a_46160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X73 VSS byte3.tinv7.I a_70320_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X74 a_98040_306# byte2.cgate0.nand0.A byte2.cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X75 a_4330_140# byte4.dff_1.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X76 a_115030_140# byte2.dff_3.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X77 VSS byte2.tinv6.I a_128640_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X78 byte4.dff_1.O byte4.dff_1.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X79 VSS a_11460_190# a_12120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X80 a_24020_1090# byte4.dff_6.CLK a_23850_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X81 byte3.dff_1.O byte3.dff_1.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X82 Do18 byte3.tinv5.ENB a_62760_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X83 VDD byte2.tinv2.I a_113520_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X84 VDD byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X85 byte4.dff_3.O byte4.dff_3.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X86 VSS a_22800_190# a_23460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X87 Do17 byte3.tinv6.EN a_66540_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X88 byte3.dff_4.O byte3.dff_4.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X89 VDD a_122160_190# a_122820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X90 a_171840_680# a_171630_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X91 VSS a_159340_140# a_159240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X92 a_163450_140# byte1.dff_5.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X93 VSS byte4.tinv5.I a_21720_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X94 VSS a_3900_190# a_4560_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X95 a_23460_1090# a_23230_140# a_22900_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X96 VDD byte2.cgate0.nand0.B byte2.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X97 VDD byte2.tinv0.I a_105960_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X98 byte1.nand.OUT WE0 a_133860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X99 VDD a_4000_140# a_3900_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X100 VSS byte4.tinv0.I a_2820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X101 VSS a_44940_190# a_45600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X102 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X103 VDD a_156720_680# a_156680_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X104 byte1.cgate0.nand0.OUT byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X105 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X106 VSS a_171840_680# a_171800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X107 VSS byte3.tinv0.I a_43860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X108 byte3.buf_RE1.O byte3.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X109 gt_re2.O gt_re2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X110 a_119600_1090# byte2.dff_4.CLK a_119430_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X111 Do27 byte4.tinv4.EN a_17940_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X112 a_115540_190# a_114600_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X113 a_158160_1092# byte1.tinv3.ENB Do4 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X114 a_41590_140# byte3.dff_0.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X115 byte2.buf_RE1.O byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X116 VDD a_163120_140# a_163020_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X117 a_126880_190# a_125940_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X118 VDD a_149160_680# a_149120_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X119 VSS byte2.cgate0.nand0.B byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X120 a_108260_190# a_107470_140# a_108090_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X121 a_27010_140# byte4.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X122 byte3.buf_RE1.O byte3.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X123 buf_ck1.O buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X124 a_121080_1092# byte2.tinv4.ENB Do11 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X125 byte1.nand.OUT WE0 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X126 a_220_140# byte4.dff_0.CLK a_450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X127 a_29280_1092# byte4.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X128 byte4.cgate0.latch0.I0.O byte4.cgate0.latch0.I0.O a_37560_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X129 a_144450_190# Di7 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X130 a_8110_140# byte4.dff_2.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X131 VDD byte3.tinv0.I a_43860_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X132 a_136020_306# byte1.cgate0.latch0.I0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X133 a_68840_190# a_68050_140# a_68670_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X134 a_155790_190# Di4 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X135 a_12680_1090# byte4.dff_3.CLK a_12510_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X136 VDD byte2.buf_RE1.I byte2.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X137 a_113520_1092# byte2.tinv2.ENB Do13 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X138 a_152730_190# byte1.dff_2.CLK a_152620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X139 VDD byte3.tinv6.I a_66540_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X140 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X141 VDD a_110820_190# a_111480_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X142 a_160500_680# a_160290_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X143 a_152110_140# byte1.dff_2.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X144 Do28 byte4.tinv3.ENB a_14160_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X145 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X146 a_107700_190# byte2.dff_1.CLK a_107140_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X147 a_168060_680# a_167850_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X148 a_27520_190# a_26580_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X149 a_49940_1090# byte3.dff_2.CLK a_49770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X150 byte2.cgate0.latch0.I0.O byte2.cgate0.nand0.B a_96420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X151 a_158160_306# byte1.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X152 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X153 VDD byte1.cgate0.nand0.A byte1.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X154 a_8010_1090# Di29 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X155 a_108260_1090# byte2.dff_1.CLK a_108090_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X156 Do5 byte1.tinv2.EN a_154380_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X157 a_8620_190# a_7680_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X158 byte1.dff_0.O byte1.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X159 VDD a_8940_680# byte4.dff_2.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X160 VSS a_4000_140# a_3900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X161 byte1.dff_3.O byte1.dff_3.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X162 a_49380_1090# a_49150_140# a_48820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X163 VSS a_45040_140# a_44940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X164 a_119640_680# a_119430_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X165 a_155560_140# byte1.dff_3.CLK a_155790_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X166 byte3.buf_RE1.O byte3.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X167 a_68280_190# byte3.dff_7.CLK a_67720_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X168 a_29280_1092# byte4.tinv7.ENB Do24 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X169 VDD a_168060_680# byte1.dff_6.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X170 VSS a_24060_680# byte4.dff_6.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X171 a_151780_140# a_152110_140# a_152010_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X172 VSS a_144120_190# a_144780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X173 VDD byte4.buf_RE0.I byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X174 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X175 VSS byte3.buf_RE0.I byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X176 VSS gt_re2.I gt_re2.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X177 a_130150_140# byte2.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X178 a_126270_190# Di9 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X179 VDD a_20280_680# a_20240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X180 VSS a_5160_680# byte4.dff_1.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X181 a_95160_1092# byte2.cgate0.latch0.I0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X182 VDD byte2.buf_RE1.I byte2.buf_RE1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X183 a_70320_306# byte3.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X184 byte2.cgate0.nand0.OUT byte2.cgate0.nand0.A a_98040_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X185 VSS a_115860_680# a_115820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X186 VDD a_41160_190# a_41820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X187 a_123210_190# byte2.dff_5.CLK a_123100_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X188 a_19680_190# byte4.dff_5.CLK a_19120_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X189 a_128640_306# byte2.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X190 VDD byte3.tinv3.I a_55200_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X191 a_66540_1092# byte3.tinv6.ENB Do17 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X192 a_81660_306# WE2 byte3.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X193 VDD a_123420_680# a_123380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X194 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X195 byte4.dff_1.O byte4.dff_1.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X196 VSS byte4.cgate0.latch0.I0.I a_37560_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X197 VDD a_63840_190# a_64500_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X198 byte1.dff_7.O byte1.dff_7.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X199 VSS a_170680_140# a_170580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X200 a_780_190# byte4.dff_0.CLK a_220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X201 VSS a_46200_680# byte3.dff_1.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X202 a_136020_306# byte1.cgate0.latch0.I0.O byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X203 a_21720_306# byte4.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X204 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X205 a_168020_190# a_167230_140# a_167850_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X206 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X207 a_8730_190# a_8110_140# a_8620_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X208 a_41490_190# Di23 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X209 a_6600_1092# byte4.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X210 byte2.buf_RE0.O byte2.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X211 a_148330_140# byte1.dff_1.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X212 a_152340_1090# a_152110_140# a_151780_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X213 byte1.buf_RE1.O byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X214 a_2820_306# byte4.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X215 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X216 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X217 a_122260_140# a_122590_140# a_122490_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X218 byte1.dff_5.O byte1.dff_5.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X219 a_7780_140# byte4.dff_2.CLK a_8010_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X220 VSS byte3.buf_RE1.I byte3.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X221 a_167850_190# a_167230_140# a_167740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X222 a_155790_1090# Di4 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X223 a_144220_140# byte1.dff_0.CLK a_144450_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X224 a_53760_680# a_53550_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X225 a_165720_1092# byte1.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X226 byte3.buf_RE0.O byte3.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X227 VSS byte2.cgate0.latch0.I0.O byte2.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X228 VSS a_114600_190# a_115260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X229 a_158160_306# byte1.tinv3.EN Do4 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X230 VDD a_156720_680# byte1.dff_3.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X231 a_149160_680# a_148950_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X232 VSS a_27840_680# a_27800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X233 a_65100_680# a_64890_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X234 VSS byte2.tinv2.I a_113520_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X235 a_62760_1092# byte3.tinv5.ENB Do18 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X236 byte2.cgate0.latch0.I0.O byte2.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X237 a_166900_140# byte1.dff_6.CLK a_167130_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X238 VSS a_171840_680# byte1.dff_7.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X239 a_148230_1090# Di6 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X240 VSS a_8940_680# a_8900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X241 a_109740_306# byte2.tinv1.EN Do14 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X242 a_138900_306# byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X243 VDD a_53760_680# a_53720_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X244 a_148840_190# a_147900_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X245 byte3.dff_0.O byte3.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X246 VSS a_49980_680# a_49940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X247 a_121080_306# byte2.tinv4.EN Do11 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X248 a_156120_190# byte1.dff_3.CLK a_155560_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X249 a_55200_1092# byte3.tinv3.ENB Do20 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X250 a_57330_190# byte3.dff_4.CLK a_57220_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X251 VSS a_144220_140# a_144120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X252 a_5120_1090# byte4.dff_1.CLK a_4950_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X253 a_171800_1090# byte1.dff_7.CLK a_171630_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X254 a_167460_190# byte1.dff_6.CLK a_166900_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X255 VDD a_60160_140# a_60060_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X256 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X257 a_68670_190# byte3.dff_7.CLK a_68560_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X258 VDD a_52500_190# a_53160_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X259 a_23740_1090# a_22800_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X260 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X261 a_17940_1092# byte4.tinv4.ENB Do27 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X262 a_70320_306# byte3.tinv7.EN Do16 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X263 VSS byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X264 Do30 byte4.tinv1.ENB a_6600_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X265 a_122260_140# byte2.dff_5.CLK a_122490_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X266 Do0 byte1.tinv7.ENB a_173280_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X267 a_164240_1090# byte1.dff_5.CLK a_164070_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X268 VDD a_15240_190# a_15900_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X269 a_20240_190# a_19450_140# a_20070_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X270 VSS CLK buf_ck0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X271 a_126880_1090# a_125940_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X272 a_128640_306# byte2.tinv6.EN Do9 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X273 VSS byte4.tinv3.I a_14160_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X274 a_96420_306# byte2.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X275 a_111760_190# a_110820_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X276 VDD byte4.tinv7.I a_29280_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X277 VDD buf_ck1.I buf_ck1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X278 a_1340_190# a_550_140# a_1170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X279 VSS byte4.tinv6.I a_25500_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X280 a_156510_190# a_155890_140# a_156400_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X281 VSS byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X282 Do2 byte1.tinv5.ENB a_165720_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X283 a_154380_1092# byte1.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X284 a_49150_140# byte3.dff_2.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X285 a_119320_1090# a_118380_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X286 VSS a_145380_680# byte1.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X287 VSS byte4.tinv1.I a_6600_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X288 a_21720_306# byte4.tinv5.EN Do26 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X289 VSS a_164280_680# a_164240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X290 VDD a_145380_680# byte1.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X291 VSS a_48720_190# a_49380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X292 VDD byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X293 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X294 VSS byte3.tinv1.I a_47640_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X295 a_53720_190# a_52930_140# a_53550_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X296 VDD a_118480_140# a_118380_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X297 a_2820_306# byte4.tinv0.EN Do31 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X298 a_75900_306# byte3.cgate0.nand0.A byte3.cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X299 VDD a_42420_680# a_42380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X300 a_119320_190# a_118380_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X301 a_20280_680# a_20070_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X302 VSS byte4.buf_RE1.I byte4.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X303 byte3.buf_RE0.O byte3.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X304 byte1.buf_RE1.O byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X305 gt_re2.O gt_re2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X306 a_137280_1092# byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X307 a_160460_1090# byte1.dff_4.CLK a_160290_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X308 a_152940_680# a_152730_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X309 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X310 VDD a_65100_680# a_65060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X311 a_123420_680# a_123210_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X312 VDD a_130980_680# byte2.dff_7.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X313 a_12400_1090# a_11460_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X314 a_12400_190# a_11460_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X315 VSS byte2.cgate0.latch0.I0.I a_95160_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X316 a_148230_190# Di6 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X317 a_122490_1090# Di10 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X318 VDD a_11560_140# a_11460_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X319 a_110920_140# byte2.dff_2.CLK a_111150_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X320 a_159570_190# Di3 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X321 Do3 byte1.tinv4.ENB a_161940_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X322 a_132420_1092# byte2.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X323 VDD a_27840_680# a_27800_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X324 a_107470_140# byte2.dff_1.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X325 a_115860_680# a_115650_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X326 VSS a_115860_680# byte2.dff_3.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X327 byte1.cgate0.latch0.I0.O byte1.cgate0.latch0.I0.O a_136020_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X328 VDD a_123420_680# byte2.dff_5.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X329 a_156510_190# byte1.dff_3.CLK a_156400_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X330 VDD byte3.buf_RE1.I byte3.buf_RE1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X331 a_159670_140# byte1.dff_4.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X332 a_45880_190# a_44940_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X333 a_53160_190# byte3.dff_3.CLK a_52600_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X334 VDD a_114700_140# a_114600_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X335 VSS byte1.tinv4.I a_161940_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X336 a_145170_190# a_144550_140# a_145060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X337 VSS a_26680_140# a_26580_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X338 byte4.buf_RE0.O byte4.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X339 Do5 byte1.tinv2.ENB a_154380_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X340 byte4.buf_RE0.O byte4.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X341 VSS byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X342 VSS byte1.tinv7.I a_173280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X343 VSS a_7780_140# a_7680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X344 byte3.buf_RE1.O byte3.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X345 a_169500_306# byte1.tinv6.EN Do1 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X346 buf_ck1.O buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X347 byte2.cgate0.nand0.A byte2.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X348 VDD a_107140_140# a_107040_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X349 a_113520_306# byte2.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X350 a_159900_1090# a_159670_140# a_159340_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X351 VSS byte3.cgate0.nand0.B byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X352 a_124860_306# byte2.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X353 a_130770_190# a_130150_140# a_130660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X354 a_155560_140# a_155890_140# a_155790_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X355 a_130050_190# Di8 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X356 VDD byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X357 a_23230_140# byte4.dff_6.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X358 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X359 a_103690_140# byte2.dff_0.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X360 Do11 byte2.tinv4.EN a_121080_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X361 VDD byte4.tinv1.I a_6600_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X362 a_52830_1090# Di20 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X363 a_37560_1092# byte4.cgate0.latch0.I0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X364 a_41260_140# byte3.dff_0.CLK a_41490_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X365 VSS a_27840_680# byte4.dff_7.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X366 VDD byte2.nand.B byte2.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X367 VDD byte2.buf_RE0.I byte2.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X368 a_152900_190# a_152110_140# a_152730_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X369 VSS a_147900_190# a_148560_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X370 a_45880_1090# a_44940_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X371 VSS a_61320_680# a_61280_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X372 a_160180_190# a_159240_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X373 VSS byte1.tinv0.I a_146820_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X374 VDD a_53760_680# byte3.dff_3.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X375 a_121080_1092# byte2.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X376 a_123210_190# a_122590_140# a_123100_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X377 VSS a_8940_680# byte4.dff_2.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X378 VDD a_16500_680# a_16460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X379 a_104520_680# a_104310_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X380 VSS byte3.buf_RE0.I byte3.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X381 VSS a_119640_680# a_119600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X382 VSS byte1.buf_RE1.I byte1.buf_RE1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X383 Do8 byte2.tinv7.ENB a_132420_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X384 a_130150_140# byte2.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X385 a_63940_140# byte3.dff_6.CLK a_64170_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X386 VDD byte3.buf_RE0.I byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X387 VDD byte1.tinv5.I a_165720_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X388 byte4.buf_RE1.O byte4.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X389 a_68560_1090# a_67620_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X390 a_68880_680# a_68670_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X391 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X392 VDD a_7680_190# a_8340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X393 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X394 buf_ck0.O CLK VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X395 VSS a_12720_680# a_12680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X396 VDD a_67720_140# a_67620_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X397 a_20070_190# byte4.dff_5.CLK a_19960_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X398 a_95160_1092# byte2.cgate0.latch0.I0.ENB byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X399 a_108300_680# a_108090_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X400 VDD byte1.tinv3.I a_158160_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X401 a_25500_306# byte4.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X402 a_45270_190# Di22 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X403 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X404 a_1170_190# byte4.dff_0.CLK a_1060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X405 Do26 byte4.tinv5.EN a_21720_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X406 VSS a_60060_190# a_60720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X407 byte2.cgate0.nand0.OUT byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X408 a_6600_306# byte4.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X409 a_42210_190# byte3.dff_0.CLK a_42100_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X410 a_148560_1090# a_148330_140# a_148000_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X411 VSS byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X412 Do16 byte3.tinv7.ENB a_70320_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X413 a_126040_140# a_126370_140# a_126270_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X414 Do31 byte4.tinv0.EN a_2820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X415 a_42420_680# a_42210_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X416 a_47640_306# byte3.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X417 byte3.cgate0.nand0.OUT byte3.cgate0.nand0.A a_75900_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X418 VDD a_49980_680# byte3.dff_2.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X419 byte4.buf_RE1.O byte4.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X420 a_57540_680# a_57330_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X421 a_58980_306# byte3.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X422 VSS byte2.tinv0.I a_105960_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X423 a_41490_1090# Di23 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X424 a_123380_190# a_122590_140# a_123210_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X425 a_6600_1092# byte4.tinv1.ENB Do30 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X426 a_53550_190# a_52930_140# a_53440_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X427 Do20 byte3.tinv3.EN a_55200_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X428 VDD WE2 byte3.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X429 byte2.inv_and.O byte2.inv_and.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X430 VDD byte2.buf_RE0.I byte2.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X431 VSS byte2.tinv3.I a_117300_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X432 VDD byte1.buf_RE1.I byte1.buf_RE1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X433 byte4.cgate0.latch0.I0.O byte4.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X434 a_51420_1092# byte3.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X435 a_56710_140# byte3.dff_4.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X436 a_65100_680# a_64890_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X437 VSS buf_ck1.I buf_ck1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X438 VSS byte2.cgate0.nand0.B a_98040_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X439 VDD a_3900_190# a_4560_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X440 VDD a_42420_680# byte3.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X441 a_113520_306# byte2.tinv2.EN Do13 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X442 a_171520_1090# a_170580_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X443 a_64170_1090# Di17 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X444 VDD byte3.buf_RE0.I byte3.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X445 a_103920_1090# a_103690_140# a_103360_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X446 a_124860_306# byte2.tinv5.EN Do10 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X447 a_170910_190# Di0 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X448 a_165720_1092# byte1.tinv5.ENB Do2 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X449 VDD byte1.tinv2.I a_154380_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X450 a_138900_306# byte1.cgate0.nand0.A byte1.cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X451 VSS byte4.tinv2.I a_10380_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X452 a_41260_140# a_41590_140# a_41490_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X453 a_57540_680# a_57330_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X454 a_64270_140# byte3.dff_6.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X455 VDD a_170680_140# a_170580_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X456 VSS a_148000_140# a_147900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X457 byte2.dff_3.O byte2.dff_3.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X458 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X459 a_52600_140# a_52930_140# a_52830_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X460 byte3.cgate0.nand0.OUT byte3.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X461 VDD a_163020_190# a_163680_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X462 VSS byte4.cgate0.nand0.B a_34860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X463 a_126600_1090# a_126370_140# a_126040_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X464 a_15340_140# byte4.dff_4.CLK a_15570_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X465 a_26910_1090# Di24 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X466 a_19960_1090# a_19020_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X467 VSS byte4.buf_RE0.I byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X468 a_122820_190# byte2.dff_5.CLK a_122260_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X469 VSS a_160500_680# a_160460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X470 a_550_140# byte4.dff_0.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X471 VDD a_27840_680# byte4.dff_7.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X472 byte2.dff_1.O byte2.dff_1.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X473 a_104200_190# a_103260_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X474 VSS a_110920_140# a_110820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X475 byte1.cgate0.latch0.I0.O byte1.cgate0.latch0.I0.O a_137280_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X476 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X477 a_173280_306# byte1.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X478 VDD a_155460_190# a_156120_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X479 a_15670_140# byte4.dff_4.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X480 a_118480_140# byte2.dff_4.CLK a_118710_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X481 a_19350_1090# Di26 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X482 VSS byte4.tinv4.I a_17940_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X483 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X484 a_109740_1092# byte2.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X485 Do1 byte1.tinv6.EN a_169500_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X486 VSS a_149160_680# byte1.dff_1.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X487 byte1.dff_4.O byte1.dff_4.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X488 a_5120_190# a_4330_140# a_4950_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X489 VSS byte4.tinv7.I a_29280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X490 VSS buf_ck1.I buf_ck1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X491 a_1060_1090# a_120_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X492 byte1.dff_7.O byte1.dff_7.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X493 a_159670_140# byte1.dff_4.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X494 VDD byte1.buf_RE0.I byte1.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X495 VSS a_60160_140# a_60060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X496 byte3.cgate0.latch0.I0.O byte3.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X497 a_25500_306# byte4.tinv6.EN Do25 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X498 a_42210_190# a_41590_140# a_42100_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X499 buf_ck0.O CLK VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X500 VSS a_168060_680# a_168020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X501 VDD byte2.tinv7.I a_132420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X502 VDD byte4.inv_and.I byte4.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X503 Do21 byte3.tinv2.ENB a_51420_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X504 a_57500_190# a_56710_140# a_57330_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X505 byte2.cgate0.latch0.I0.O byte2.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X506 VSS a_118480_140# a_118380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X507 VDD a_152940_680# a_152900_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X508 a_6600_306# byte4.tinv1.EN Do30 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X509 VDD RE gt_re0.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X510 a_160180_1090# a_159240_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X511 VSS a_129820_140# a_129720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X512 a_47640_306# byte3.tinv1.EN Do22 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X513 a_115820_1090# byte2.dff_3.CLK a_115650_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X514 a_12120_1090# a_11890_140# a_11560_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X515 VSS a_112080_680# byte2.dff_2.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X516 a_154380_1092# byte1.tinv2.ENB Do5 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X517 a_146820_306# byte1.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X518 VSS a_130980_680# a_130940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X519 VSS a_11560_140# a_11460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X520 byte4.dff_6.O byte4.dff_6.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X521 VSS byte4.buf_RE1.I byte4.buf_RE1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X522 a_58980_306# byte3.tinv4.EN Do19 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X523 byte2.dff_0.O byte2.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X524 a_156720_680# a_156510_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X525 a_56940_1090# a_56710_140# a_56380_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X526 byte3.cgate0.nand0.A byte3.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X527 VDD a_145380_680# a_145340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X528 VSS a_22900_140# a_22800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X529 a_15570_1090# Di27 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X530 a_16180_190# a_15240_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X531 a_27630_190# a_27010_140# a_27520_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X532 byte3.dff_7.O byte3.dff_7.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X533 a_105960_1092# byte2.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X534 a_115260_1090# a_115030_140# a_114700_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X535 Do12 byte2.tinv3.ENB a_117300_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X536 a_25500_1092# byte4.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X537 byte2.buf_RE0.O byte2.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X538 VDD a_16500_680# byte4.dff_4.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X539 VSS a_61320_680# byte3.dff_5.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X540 a_56940_190# byte3.dff_4.CLK a_56380_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X541 VDD a_168060_680# a_168020_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X542 byte1.cgate0.nand0.A byte1.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X543 a_26680_140# byte4.dff_7.CLK a_26910_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X544 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X545 a_109740_1092# byte2.tinv1.ENB Do14 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X546 a_163450_140# byte1.dff_5.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X547 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X548 a_450_1090# Di31 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X549 a_49660_190# a_48720_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X550 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X551 a_114930_190# Di12 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X552 VDD byte3.tinv5.I a_62760_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X553 VDD a_130980_680# a_130940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X554 VSS a_12720_680# byte4.dff_3.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X555 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X556 VDD byte2.tinv4.I a_121080_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X557 a_132420_1092# byte2.tinv7.ENB Do8 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X558 buf_ck1.O buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X559 a_173280_306# byte1.tinv7.EN Do0 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X560 VSS a_129720_190# a_130380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X561 VDD byte4.buf_RE1.I byte4.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X562 byte3.buf_RE0.O byte3.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X563 gt_re1.O gt_re1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X564 VSS a_104520_680# a_104480_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X565 VDD a_129720_190# a_130380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X566 a_171010_140# byte1.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X567 a_104480_1090# byte2.dff_0.CLK a_104310_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X568 a_117300_306# byte2.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X569 VDD byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X570 buf_ck1.O buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X571 VDD a_5160_680# byte4.dff_1.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X572 a_68840_1090# byte3.dff_7.CLK a_68670_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X573 Do13 byte2.tinv2.EN a_113520_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X574 a_159340_140# a_159670_140# a_159570_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X575 a_20280_680# a_20070_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X576 a_45600_1090# a_45370_140# a_45040_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X577 VSS byte3.inv_and.I byte3.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X578 a_171240_190# byte1.dff_7.CLK a_170680_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X579 a_127160_1090# byte2.dff_6.CLK a_126990_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X580 Do10 byte2.tinv5.EN a_124860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X581 a_145340_190# a_144550_140# a_145170_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X582 byte1.cgate0.nand0.OUT byte1.cgate0.nand0.A a_138900_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X583 a_16290_190# a_15670_140# a_16180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X584 byte3.dff_4.O byte3.dff_4.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X585 VDD byte2.cgate0.nand0.A byte2.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X586 Do15 byte2.tinv0.ENB a_105960_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X587 VSS buf_sel1.I buf_sel1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X588 byte2.dff_3.O byte2.dff_3.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X589 a_1380_680# a_1170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X590 a_14160_1092# byte4.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X591 a_10380_306# byte4.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X592 Do25 byte4.tinv6.ENB a_25500_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X593 a_156680_190# a_155890_140# a_156510_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X594 VSS a_65100_680# a_65060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X595 a_34860_306# byte4.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X596 a_58980_1092# byte3.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X597 a_68280_1090# a_68050_140# a_67720_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X598 a_26910_190# Di24 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X599 VSS a_103260_190# a_103920_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X600 a_146820_306# byte1.tinv0.EN Do7 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X601 a_133860_306# byte1.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X602 byte4.buf_RE0.O byte4.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X603 buf_sel0.O buf_sel0.I VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=1.02p ps=4.6u w=1.7u l=300n
X604 a_110920_140# a_111250_140# a_111150_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X605 Do9 byte2.tinv6.ENB a_128640_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X606 byte1.buf_RE0.O byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X607 a_23850_190# byte4.dff_6.CLK a_23740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X608 a_148840_1090# a_147900_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X609 a_8010_190# Di29 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X610 byte3.dff_6.O byte3.dff_6.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X611 VDD byte4.cgate0.nand0.B byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X612 a_43860_306# byte3.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X613 VDD byte3.tinv2.I a_51420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X614 a_49050_190# Di21 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X615 VDD byte2.inv_and.I byte2.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X616 a_4950_190# byte4.dff_1.CLK a_4840_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X617 VSS a_16500_680# a_16460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X618 VSS byte4.nand.B a_40620_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X619 VSS byte2.buf_RE1.I byte2.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X620 VDD a_60060_190# a_60720_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X621 buf_ck1.O buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X622 byte4.dff_0.O byte4.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X623 a_29280_306# byte4.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X624 VSS a_160500_680# byte1.dff_4.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X625 gt_re2.O gt_re2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X626 VDD a_112080_680# a_112040_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X627 a_4950_190# a_4330_140# a_4840_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X628 Do25 byte4.tinv6.EN a_25500_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X629 VSS a_63840_190# a_64500_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X630 a_2820_1092# byte4.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X631 byte4.dff_4.O byte4.dff_4.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X632 VSS byte3.tinv5.I a_62760_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X633 VDD byte3.cgate0.nand0.B byte3.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X634 VDD byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X635 a_49150_140# byte3.dff_2.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X636 buf_sel0.O buf_sel0.I VSS VSS nfet_03v3 ad=510f pd=2.9u as=510f ps=2.9u w=850n l=300n
X637 Do30 byte4.tinv1.EN a_6600_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X638 byte4.dff_7.O byte4.dff_7.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X639 a_57500_1090# byte3.dff_4.CLK a_57330_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X640 a_107470_140# byte2.dff_1.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X641 byte1.dff_4.O byte1.dff_4.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X642 a_60490_140# byte3.dff_5.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X643 a_4000_140# byte4.dff_1.CLK a_4230_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X644 VSS byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X645 a_118810_140# byte2.dff_4.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X646 a_152010_1090# Di5 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X647 byte4.dff_2.O byte4.dff_2.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X648 VDD byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X649 a_171240_1090# a_171010_140# a_170680_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X650 a_161940_1092# byte1.tinv4.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X651 a_127160_190# a_126370_140# a_126990_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X652 a_8940_680# a_8730_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X653 VSS a_15240_190# a_15900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X654 byte4.buf_RE1.O byte4.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X655 Do19 byte3.tinv4.EN a_58980_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X656 a_145380_680# a_145170_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X657 a_22900_140# a_23230_140# a_23130_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X658 a_49770_190# a_49150_140# a_49660_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X659 VDD a_152940_680# byte1.dff_2.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X660 Do19 byte3.tinv4.ENB a_58980_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X661 VDD byte3.buf_RE1.I byte3.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X662 VDD byte2.tinv1.I a_109740_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X663 a_117300_306# byte2.tinv3.EN Do12 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X664 a_163350_190# Di2 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X665 gt_re0.OUT gt_re0.A a_84900_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X666 a_4000_140# a_4330_140# a_4230_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X667 VSS byte2.buf_RE0.I byte2.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X668 a_163120_140# byte1.dff_5.CLK a_163350_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X669 a_144450_1090# Di7 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X670 byte1.buf_RE0.O byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X671 a_11890_140# byte4.dff_3.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X672 VDD buf_sel1.I buf_sel1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X673 a_168060_680# a_167850_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X674 a_45040_140# a_45370_140# a_45270_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X675 a_68050_140# byte3.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X676 a_19680_1090# a_19450_140# a_19120_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X677 a_51420_1092# byte3.tinv2.ENB Do21 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X678 VDD CLK buf_ck0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X679 VDD byte2.cgate0.nand0.B byte2.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X680 byte2.buf_RE1.O byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X681 a_171630_190# byte1.dff_7.CLK a_171520_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X682 a_1340_1090# byte4.dff_0.CLK a_1170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X683 a_10380_306# byte4.tinv2.EN Do29 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X684 a_56380_140# a_56710_140# a_56610_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X685 VDD a_166900_140# a_166800_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X686 a_167130_1090# Di1 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X687 a_61000_190# a_60060_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X688 VSS a_103360_140# a_103260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X689 a_42380_190# a_41590_140# a_42210_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X690 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X691 VSS byte4.cgate0.latch0.I0.O byte4.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X692 a_126600_190# byte2.dff_6.CLK a_126040_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X693 VSS a_114700_140# a_114600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X694 VSS byte1.inv_and.I byte1.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X695 VDD a_159340_140# a_159240_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X696 Do31 byte4.tinv0.ENB a_2820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X697 VDD byte4.cgate0.nand0.A byte4.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X698 a_43860_306# byte3.tinv0.EN Do23 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X699 VDD byte3.cgate0.latch0.I0.O byte3.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X700 byte1.dff_5.O byte1.dff_5.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X701 a_46160_1090# byte3.dff_1.CLK a_45990_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X702 gt_re2.O gt_re2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X703 byte1.dff_1.O byte1.dff_1.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X704 VDD byte4.tinv6.I a_25500_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X705 byte4.cgate0.latch0.I0.O byte4.cgate0.latch0.I0.ENB a_37560_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X706 a_152730_190# a_152110_140# a_152620_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X707 a_155890_140# byte1.dff_3.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X708 a_150600_1092# byte1.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X709 VDD byte1.cgate0.latch0.I0.O byte1.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X710 VSS byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X711 a_115540_1090# a_114600_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X712 VSS a_151680_190# a_152340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X713 Do22 byte3.tinv1.ENB a_47640_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X714 a_41820_190# byte3.dff_0.CLK a_41260_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X715 VSS a_163020_190# a_163680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X716 VDD byte4.tinv4.I a_17940_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X717 buf_sel1.O buf_sel1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X718 VSS a_104520_680# byte2.dff_0.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X719 a_170680_140# a_171010_140# a_170910_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X720 a_37560_306# byte4.cgate0.latch0.I0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X721 a_173280_1092# byte1.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X722 a_151780_140# byte1.dff_2.CLK a_152010_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X723 a_145170_190# byte1.dff_0.CLK a_145060_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X724 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X725 VDD a_107040_190# a_107700_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X726 a_156720_680# a_156510_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X727 a_148330_140# byte1.dff_1.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X728 VDD a_26580_190# a_27240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X729 a_27240_190# byte4.dff_7.CLK a_26680_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X730 VDD a_164280_680# byte1.dff_5.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X731 a_780_1090# a_550_140# a_220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X732 VSS a_15340_140# a_15240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X733 VDD buf_ck1.I buf_ck1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X734 VDD byte2.cgate0.latch0.I0.I a_95160_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X735 Do7 byte1.tinv0.EN a_146820_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X736 a_8340_190# byte4.dff_2.CLK a_7780_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X737 VSS byte4.buf_RE0.I byte4.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X738 a_136020_1092# byte1.cgate0.latch0.I0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X739 VDD a_61320_680# a_61280_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X740 VDD gt_re1.I gt_re1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X741 Do4 byte1.tinv3.EN a_158160_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X742 a_112080_680# a_111870_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X743 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X744 byte1.buf_RE0.O byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X745 byte2.buf_RE1.O byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X746 a_123420_680# a_123210_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X747 VDD a_148000_140# a_147900_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X748 a_40620_306# WE3 byte4.nand.OUT VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X749 VSS a_48820_140# a_48720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X750 a_60390_190# Di18 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X751 a_78240_1092# byte3.cgate0.latch0.I0.O byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X752 a_111760_1090# a_110820_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X753 a_112080_680# a_111870_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X754 a_167230_140# byte1.dff_6.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X755 a_144220_140# a_144550_140# a_144450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X756 VDD a_119640_680# byte2.dff_4.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X757 a_118710_190# Di11 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X758 byte3.inv_and.O byte3.inv_and.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X759 a_105960_1092# byte2.tinv0.ENB Do15 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X760 a_25500_1092# byte4.tinv6.ENB Do25 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X761 VDD a_110920_140# a_110820_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X762 Do14 byte2.tinv1.EN a_109740_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X763 a_111150_1090# Di13 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X764 a_115650_190# byte2.dff_3.CLK a_115540_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X765 a_129820_140# byte2.dff_7.CLK a_130050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X766 Do6 byte1.tinv1.ENB a_150600_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X767 VDD byte1.cgate0.nand0.B byte1.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X768 VSS a_16500_680# byte4.dff_4.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X769 VDD a_22800_190# a_23460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X770 VSS byte4.cgate0.nand0.A a_37200_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X771 a_104200_1090# a_103260_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X772 a_126370_140# byte2.dff_6.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X773 a_126990_190# byte2.dff_6.CLK a_126880_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X774 a_11790_190# Di28 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X775 byte4.cgate0.inv1.O byte4.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X776 VSS a_108300_680# a_108260_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X777 VDD byte1.buf_RE0.I byte1.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X778 byte4.dff_2.O byte4.dff_2.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X779 Do16 byte3.tinv7.EN a_70320_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X780 a_164070_190# a_163450_140# a_163960_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X781 VSS byte2.tinv7.I a_132420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X782 VDD a_103360_140# a_103260_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X783 VDD a_119640_680# a_119600_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X784 byte2.dff_1.O byte2.dff_1.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X785 a_167740_190# a_166800_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X786 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X787 a_24060_680# a_23850_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X788 byte3.dff_5.O byte3.dff_5.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X789 VSS a_68880_680# a_68840_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X790 VSS a_163120_140# a_163020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X791 a_149120_190# a_148330_140# a_148950_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X792 byte2.buf_RE0.O byte2.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X793 VDD a_126040_140# a_125940_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X794 Do9 byte2.tinv6.EN a_128640_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X795 a_14160_306# byte4.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X796 a_19450_140# byte4.dff_5.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X797 byte4.buf_RE0.O byte4.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X798 VDD gt_re2.I gt_re2.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X799 byte1.cgate0.latch0.I0.O byte1.cgate0.latch0.I0.ENB a_136020_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X800 VDD byte4.tinv0.I a_2820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X801 a_5160_680# a_4950_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X802 a_19350_190# Di26 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X803 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X804 byte2.nand.OUT WE1 a_93000_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X805 Do29 byte4.tinv2.EN a_10380_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X806 VSS byte4.cgate0.nand0.B byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X807 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X808 VSS a_107040_190# a_107700_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X809 a_450_190# Di31 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X810 VDD a_12720_680# a_12680_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X811 byte4.cgate0.nand0.A byte4.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X812 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X813 a_112040_190# a_111250_140# a_111870_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X814 a_114700_140# a_115030_140# a_114930_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X815 a_122590_140# byte2.dff_5.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X816 byte4.dff_3.O byte4.dff_3.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X817 a_27630_190# byte4.dff_7.CLK a_27520_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X818 byte1.inv_and.O byte1.inv_and.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X819 a_60160_140# byte3.dff_5.CLK a_60390_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X820 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X821 a_130660_190# a_129720_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X822 a_14160_1092# byte4.tinv3.ENB Do28 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X823 a_64780_1090# a_63840_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X824 a_103690_140# byte2.dff_0.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X825 a_8730_190# byte4.dff_2.CLK a_8620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X826 Do23 byte3.tinv0.EN a_43860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X827 a_58980_1092# byte3.tinv4.ENB Do19 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X828 a_115030_140# byte2.dff_3.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X829 a_8900_1090# byte4.dff_2.CLK a_8730_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X830 VDD a_63940_140# a_63840_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X831 buf_sel1.O buf_sel1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X832 VDD byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X833 VSS byte2.buf_RE1.I byte2.buf_RE1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X834 VSS a_164280_680# byte1.dff_5.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X835 a_159900_190# byte1.dff_4.CLK a_159340_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X836 VDD byte1.buf_RE0.I byte1.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X837 VDD a_49980_680# a_49940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X838 a_57220_1090# a_56280_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X839 VSS a_67620_190# a_68280_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X840 VDD byte2.buf_RE1.I byte2.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X841 VSS byte3.tinv6.I a_66540_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X842 a_95160_306# byte2.cgate0.latch0.I0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X843 VDD a_108300_680# a_108260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X844 a_168020_1090# byte1.dff_6.CLK a_167850_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X845 a_144780_1090# a_144550_140# a_144220_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X846 VDD a_56380_140# a_56280_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X847 VDD a_48720_190# a_49380_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X848 VSS buf_sel1.I buf_sel1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X849 a_161940_306# byte1.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X850 byte1.dff_3.O byte1.dff_3.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X851 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X852 VDD byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X853 VDD gt_re2.I gt_re2.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X854 a_111480_190# byte2.dff_2.CLK a_110920_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X855 a_171840_680# a_171630_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X856 VSS a_19020_190# a_19680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X857 a_34860_306# byte4.cgate0.nand0.A byte4.cgate0.nand0.OUT VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X858 a_130050_1090# Di8 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X859 a_167460_1090# a_167230_140# a_166900_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X860 a_2820_1092# byte4.tinv0.ENB Do31 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X861 a_24020_190# a_23230_140# a_23850_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X862 a_26680_140# a_27010_140# a_26910_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X863 VSS byte3.buf_RE1.I byte3.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X864 a_52930_140# byte3.dff_3.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X865 a_61320_680# a_61110_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X866 a_167130_190# Di1 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X867 VSS a_120_190# a_780_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X868 a_7780_140# a_8110_140# a_8010_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X869 a_37560_1092# byte4.cgate0.latch0.I0.ENB byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X870 byte1.dff_1.O byte1.dff_1.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X871 VSS byte1.buf_RE0.I byte1.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X872 a_48820_140# a_49150_140# a_49050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X873 a_53440_190# a_52500_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X874 a_60390_1090# Di18 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X875 a_161940_1092# byte1.tinv4.ENB Do3 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X876 VDD byte1.tinv1.I a_150600_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X877 a_45370_140# byte3.dff_1.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X878 a_70320_1092# byte3.tinv7.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X879 a_14160_306# byte4.tinv3.EN Do28 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X880 a_53760_680# a_53550_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X881 VDD a_61320_680# byte3.dff_5.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X882 a_64780_190# a_63840_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X883 VSS a_107140_140# a_107040_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X884 a_46160_190# a_45370_140# a_45990_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X885 VDD a_52600_140# a_52500_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X886 a_11560_140# byte4.dff_3.CLK a_11790_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X887 a_122820_1090# a_122590_140# a_122260_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X888 VDD byte1.tinv7.I a_173280_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X889 a_145380_680# a_145170_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X890 VDD byte1.buf_RE1.I byte1.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X891 a_68050_140# byte3.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X892 VDD a_24060_680# byte4.dff_6.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X893 a_37200_306# byte4.cgate0.nand0.B byte4.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X894 a_12120_190# byte4.dff_3.CLK a_11560_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X895 buf_ck1.O buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X896 byte3.buf_RE0.O byte3.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X897 VDD a_151680_190# a_152340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X898 VSS byte1.cgate0.nand0.B byte1.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X899 VSS byte4.cgate0.nand0.OUT byte4.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X900 byte1.dff_6.O byte1.dff_6.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X901 a_156680_1090# byte1.dff_3.CLK a_156510_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X902 VDD a_45040_140# a_44940_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X903 byte2.cgate0.nand0.OUT byte2.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X904 a_132420_306# byte2.tinv7.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X905 a_23460_190# byte4.dff_6.CLK a_22900_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X906 byte2.dff_6.O byte2.dff_6.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X907 byte1.buf_RE1.O byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X908 a_148950_190# byte1.dff_1.CLK a_148840_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X909 a_4560_190# byte4.dff_1.CLK a_4000_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X910 a_118710_1090# Di11 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X911 VSS a_155460_190# a_156120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X912 a_149120_1090# byte1.dff_1.CLK a_148950_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X913 a_45600_190# byte3.dff_1.CLK a_45040_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X914 a_107140_140# byte2.dff_1.CLK a_107370_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X915 a_128640_1092# byte2.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X916 Do4 byte1.tinv3.ENB a_158160_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X917 VSS byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X918 byte2.dff_7.O byte2.dff_7.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X919 a_41590_140# byte3.dff_0.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X920 VDD byte3.cgate0.nand0.A a_78240_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X921 VSS a_108300_680# byte2.dff_1.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X922 VSS a_166800_190# a_167460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X923 a_171800_190# a_171010_140# a_171630_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X924 a_95160_306# byte2.cgate0.latch0.I0.O byte2.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X925 VSS byte1.tinv5.I a_165720_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X926 VDD byte4.cgate0.latch0.I0.I a_37560_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X927 a_152110_140# byte1.dff_2.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X928 a_78600_306# byte3.cgate0.latch0.I0.O byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X929 a_103590_190# Di15 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X930 a_112040_1090# byte2.dff_2.CLK a_111870_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X931 VSS a_19120_140# a_19020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X932 byte4.cgate0.latch0.I0.O byte4.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X933 a_61110_190# a_60490_140# a_61000_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X934 a_161940_306# byte1.tinv4.EN Do3 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X935 a_150600_1092# byte1.tinv1.ENB Do6 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X936 byte1.cgate0.latch0.I0.O byte1.cgate0.nand0.B a_137280_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X937 byte1.buf_RE0.O byte1.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X938 VDD a_5160_680# a_5120_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X939 byte4.dff_5.O byte4.dff_5.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X940 VSS a_20280_680# a_20240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X941 VDD a_171840_680# a_171800_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X942 a_111870_190# byte2.dff_2.CLK a_111760_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X943 VSS a_220_140# a_120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X944 a_11790_1090# Di28 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X945 a_23850_190# a_23230_140# a_23740_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X946 a_111480_1090# a_111250_140# a_110920_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X947 a_115860_680# a_115650_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X948 a_173280_1092# byte1.tinv7.ENB Do0 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X949 VSS a_1380_680# a_1340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X950 a_21720_1092# byte4.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X951 a_98040_306# byte2.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X952 VDD a_12720_680# byte4.dff_3.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X953 byte2.dff_5.O byte2.dff_5.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X954 a_127200_680# a_126990_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X955 buf_ck1.O buf_ck1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X956 a_64170_190# Di17 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X957 VDD a_164280_680# a_164240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X958 a_126990_190# a_126370_140# a_126880_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X959 a_148000_140# a_148330_140# a_148230_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X960 a_22900_140# byte4.dff_6.CLK a_23130_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X961 VSS a_53760_680# a_53720_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X962 gt_re2.O gt_re2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X963 a_124860_1092# byte2.tinv5.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X964 a_152620_190# a_151680_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X965 a_136020_1092# byte1.cgate0.latch0.I0.ENB byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X966 a_61110_190# byte3.dff_5.CLK a_61000_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X967 a_108300_680# a_108090_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X968 a_27840_680# a_27630_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X969 a_49050_1090# Di21 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X970 a_66540_306# byte3.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X971 byte2.dff_0.O byte2.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X972 a_119430_190# byte2.dff_4.CLK a_119320_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X973 a_163960_190# a_163020_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X974 a_107370_1090# Di14 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X975 a_117300_1092# byte2.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X976 a_119430_190# a_118810_140# a_119320_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X977 a_15570_190# Di27 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X978 VSS byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X979 VDD a_108300_680# byte2.dff_1.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X980 a_42420_680# a_42210_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X981 byte3.nand.OUT byte3.nand.B VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X982 a_12510_190# byte4.dff_3.CLK a_12400_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X983 byte2.cgate0.inv1.O byte2.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X984 a_132420_306# byte2.tinv7.EN Do8 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X985 VDD a_19120_140# a_19020_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X986 a_20240_1090# byte4.dff_5.CLK a_20070_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X987 a_17940_306# byte4.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X988 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X989 a_27840_680# a_27630_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X990 a_41820_1090# a_41590_140# a_41260_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X991 a_60160_140# a_60490_140# a_60390_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X992 VDD buf_sel1.I buf_sel1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X993 VDD a_160500_680# a_160460_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X994 a_123380_1090# byte2.dff_5.CLK a_123210_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X995 byte1.buf_RE0.O byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X996 a_12510_190# a_11890_140# a_12400_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X997 a_8940_680# a_8730_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X998 byte3.dff_3.O byte3.dff_3.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X999 byte2.buf_RE1.O byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1000 a_144780_190# byte1.dff_0.CLK a_144220_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1001 a_10380_1092# byte4.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1002 Do26 byte4.tinv5.ENB a_21720_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1003 a_45990_190# byte3.dff_1.CLK a_45880_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1004 VSS a_52500_190# a_53160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1005 VSS byte3.tinv2.I a_51420_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1006 a_64500_1090# a_64270_140# a_63940_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1007 a_115820_190# a_115030_140# a_115650_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1008 VSS byte2.tinv1.I a_109740_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1009 a_123100_190# a_122160_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1010 a_8620_1090# a_7680_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1011 a_11560_140# a_11890_140# a_11790_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1012 byte3.dff_1.O byte3.dff_1.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1013 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1014 VSS byte3.cgate0.nand0.B a_75900_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1015 Do10 byte2.tinv5.ENB a_124860_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1016 VSS byte1.cgate0.latch0.I0.O byte1.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1017 VDD byte4.buf_RE0.I byte4.buf_RE0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1018 VSS a_168060_680# byte1.dff_6.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1019 a_16500_680# a_16290_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1020 a_56380_140# byte3.dff_4.CLK a_56610_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1021 VSS byte3.buf_RE0.I byte3.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1022 byte1.cgate0.latch0.I0.O byte1.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1023 byte4.cgate0.nand0.OUT byte4.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1024 a_47640_1092# byte3.tinv1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1025 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1026 VDD a_7780_140# a_7680_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1027 Do22 byte3.tinv1.EN a_47640_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1028 VDD a_68880_680# byte3.dff_7.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1029 a_108090_190# a_107470_140# a_107980_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1030 a_167740_1090# a_166800_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1031 VSS byte1.buf_RE1.I byte1.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1032 a_48820_140# byte3.dff_2.CLK a_49050_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1033 VDD byte3.tinv7.I a_70320_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1034 VSS a_119640_680# byte2.dff_4.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1035 byte1.cgate0.inv1.O byte1.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1036 a_160290_190# byte1.dff_4.CLK a_160180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1037 VDD a_159240_190# a_159900_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1038 VSS a_152940_680# a_152900_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1039 VDD a_220_140# a_120_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1040 byte4.buf_RE1.O byte4.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1041 a_66540_306# byte3.tinv6.EN Do17 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1042 a_53720_1090# byte3.dff_3.CLK a_53550_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1043 a_165720_306# byte1.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1044 VSS a_130980_680# byte2.dff_7.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1045 byte2.nand.OUT WE1 VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1046 byte2.buf_RE0.O byte2.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1047 byte3.cgate0.latch0.I0.O byte3.cgate0.latch0.I0.O a_78600_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1048 byte1.buf_RE1.O byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1049 a_107980_190# a_107040_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1050 a_115260_190# byte2.dff_3.CLK a_114700_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1051 byte3.dff_0.O byte3.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1052 a_27800_190# a_27010_140# a_27630_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1053 a_137280_306# byte1.cgate0.nand0.A VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1054 VDD byte1.nand.B byte1.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1055 a_5160_680# a_4950_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1056 Do29 byte4.tinv2.ENB a_10380_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1057 Do0 byte1.tinv7.EN a_173280_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1058 a_45990_190# a_45370_140# a_45880_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1059 a_8900_190# a_8110_140# a_8730_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1060 a_43860_1092# byte3.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1061 a_53160_1090# a_52930_140# a_52600_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1062 Do20 byte3.tinv3.ENB a_55200_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1063 a_4230_1090# Di30 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1064 a_17940_306# byte4.tinv4.EN Do27 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1065 a_170910_1090# Di0 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1066 a_49940_190# a_49150_140# a_49770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1067 VSS a_63940_140# a_63840_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1068 VSS buf_ck1.I buf_ck1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1069 a_163960_1090# a_163020_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1070 a_57220_190# a_56280_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1071 byte3.cgate0.nand0.OUT byte3.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1072 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1073 a_164280_680# a_164070_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1074 a_68670_190# a_68050_140# a_68560_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1075 VDD a_171840_680# byte1.dff_7.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1076 VSS byte1.buf_RE0.I byte1.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1077 a_15900_1090# a_15670_140# a_15340_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1078 byte4.cgate0.nand0.A byte4.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1079 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1080 a_68560_190# a_67620_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1081 byte3.inv_and.O byte3.inv_and.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1082 VDD byte2.tinv6.I a_128640_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1083 byte4.dff_7.O byte4.dff_7.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1084 a_163350_1090# Di2 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1085 a_156400_1090# a_155460_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1086 a_149160_680# a_148950_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1087 VSS a_112080_680# a_112040_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1088 VSS byte1.tinv1.I a_150600_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1089 a_70320_1092# byte3.tinv7.ENB Do16 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1090 VSS a_123420_680# a_123380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1091 VDD a_155560_140# a_155460_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1092 a_19960_190# a_19020_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1093 byte4.buf_RE1.O byte4.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1094 VSS a_53760_680# byte3.dff_3.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1095 VDD byte3.buf_RE0.I byte3.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1096 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1097 VDD a_147900_190# a_148560_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1098 VSS byte1.cgate0.latch0.I0.I a_136020_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1099 VDD byte4.tinv5.I a_21720_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1100 a_42380_1090# byte3.dff_0.CLK a_42210_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1101 Do8 byte2.tinv7.EN a_132420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1102 VSS a_65100_680# byte3.dff_6.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1103 VSS byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1104 a_164240_190# a_163450_140# a_164070_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1105 byte1.inv_and.O byte1.inv_and.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1106 VDD a_1380_680# byte4.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1107 a_49380_190# byte3.dff_2.CLK a_48820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1108 VDD buf_ck1.I buf_ck1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1109 a_96420_1092# byte2.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1110 VSS byte1.tinv3.I a_158160_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1111 a_65060_1090# byte3.dff_6.CLK a_64890_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1112 Do23 byte3.tinv0.ENB a_43860_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1113 VDD gt_re2.I gt_re2.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1114 VSS byte1.tinv6.I a_169500_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1115 VDD byte4.tinv3.I a_14160_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1116 a_171630_190# a_171010_140# a_171520_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1117 a_8110_140# byte4.dff_2.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1118 a_107370_190# Di14 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1119 a_165720_306# byte1.tinv5.EN Do2 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1120 VDD a_103260_190# a_103920_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1121 VSS a_122160_190# a_122820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1122 a_152940_680# a_152730_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1123 a_129820_140# a_130150_140# a_130050_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1124 a_144550_140# byte1.dff_0.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1125 a_51420_306# byte3.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1126 VSS byte3.cgate0.latch0.I0.I a_78600_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1127 a_104310_190# byte2.dff_0.CLK a_104200_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1128 VDD a_160500_680# byte1.dff_4.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1129 a_27800_1090# byte4.dff_7.CLK a_27630_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1130 Do17 byte3.tinv6.ENB a_66540_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1131 a_109740_306# byte2.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1132 VDD byte2.tinv3.I a_117300_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1133 a_128640_1092# byte2.tinv6.ENB Do9 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1134 VSS a_24060_680# a_24020_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1135 a_62760_306# byte3.tinv5.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1136 a_75900_306# byte3.cgate0.nand0.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1137 byte1.cgate0.nand0.A byte1.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1138 a_67950_190# Di16 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1139 a_170680_140# byte1.dff_7.CLK a_170910_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1140 VSS byte2.tinv4.I a_121080_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1141 VDD a_125940_190# a_126600_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1142 a_167230_140# byte1.dff_6.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1143 a_145060_1090# a_144120_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1144 VSS a_5160_680# a_5120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1145 byte3.dff_2.O byte3.dff_2.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1146 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1147 Do24 byte4.tinv7.ENB a_29280_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1148 Do12 byte2.tinv3.EN a_117300_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1149 VSS a_151780_140# a_151680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1150 a_84900_306# RE VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1151 VDD a_144220_140# a_144120_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1152 VSS byte4.buf_RE1.I byte4.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1153 a_156400_190# a_155460_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1154 VSS a_57540_680# a_57500_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1155 VSS byte3.nand.B a_81660_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1156 VDD a_118380_190# a_119040_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1157 byte1.buf_RE1.O byte1.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1158 a_12720_680# a_12510_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1159 VDD byte4.tinv2.I a_10380_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1160 a_1170_190# a_550_140# a_1060_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1161 a_21720_1092# byte4.tinv5.ENB Do26 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1162 a_103360_140# a_103690_140# a_103590_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1163 VSS byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1164 a_126370_140# byte2.dff_6.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1165 gt_re0.OUT gt_re0.A VDD VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1166 a_130660_1090# a_129720_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1167 byte1.cgate0.latch0.I0.O byte1.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1168 a_130980_680# a_130770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1169 byte3.dff_7.O byte3.dff_7.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1170 a_124860_1092# byte2.tinv5.ENB Do10 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1171 a_16290_190# byte4.dff_4.CLK a_16180_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1172 a_46200_680# a_45990_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1173 a_160290_190# a_159670_140# a_160180_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1174 a_19450_140# byte4.dff_5.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1175 VSS byte3.cgate0.nand0.OUT byte3.cgate0.inv1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1176 Do1 byte1.tinv6.ENB a_169500_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1177 VDD byte4.cgate0.nand0.B byte4.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1178 VDD byte3.tinv1.I a_47640_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1179 VDD a_115860_680# a_115820_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1180 a_123100_1090# a_122160_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1181 VSS a_152940_680# byte1.dff_2.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1182 VDD a_11460_190# a_12120_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1183 VSS gt_re2.I gt_re2.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1184 a_550_140# byte4.dff_0.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1185 a_16460_1090# byte4.dff_4.CLK a_16290_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1186 VSS a_56280_190# a_56940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1187 a_63940_140# a_64270_140# a_64170_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1188 a_117300_1092# byte2.tinv3.ENB Do12 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1189 VDD a_56280_190# a_56940_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1190 byte3.cgate0.latch0.I0.O byte3.cgate0.nand0.B VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1191 Do24 byte4.tinv7.EN a_29280_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1192 buf_ck1.O buf_ck1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1193 VDD a_122260_140# a_122160_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1194 a_29280_306# byte4.tinv7.EN Do24 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1195 a_49770_190# byte3.dff_2.CLK a_49660_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1196 VDD a_114600_190# a_115260_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1197 a_148560_190# byte1.dff_1.CLK a_148000_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1198 a_8340_1090# a_8110_140# a_7780_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1199 a_52930_140# byte3.dff_3.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1200 VSS a_122260_140# a_122160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1201 byte1.buf_RE0.O byte1.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1202 Do27 byte4.tinv4.ENB a_17940_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1203 VDD byte4.buf_RE1.I byte4.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1204 VSS byte3.tinv3.I a_55200_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1205 a_61280_190# a_60490_140# a_61110_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1206 VDD byte1.cgate0.nand0.OUT byte1.cgate0.inv1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1207 a_119600_190# a_118810_140# a_119430_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1208 VDD byte1.buf_RE1.I byte1.buf_RE1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1209 a_15340_140# a_15670_140# a_15570_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1210 a_51420_306# byte3.tinv2.EN Do21 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1211 VDD byte2.buf_RE0.I byte2.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1212 a_150600_306# byte1.tinv1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1213 a_62760_306# byte3.tinv5.EN Do18 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1214 byte2.cgate0.latch0.I0.O byte2.cgate0.latch0.I0.ENB a_95160_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1215 VSS byte3.cgate0.latch0.I0.O byte3.cgate0.nand0.A VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1216 a_160500_680# a_160290_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1217 VSS byte1.cgate0.nand0.B a_138900_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1218 a_10380_1092# byte4.tinv2.ENB Do29 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1219 a_61000_1090# a_60060_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1220 VDD a_149160_680# byte1.dff_1.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1221 a_12680_190# a_11890_140# a_12510_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1222 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1223 a_111250_140# byte2.dff_2.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1224 a_119640_680# a_119430_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1225 VSS a_170580_190# a_171240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1226 a_159340_140# byte1.dff_4.CLK a_159570_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1227 VDD byte3.cgate0.nand0.A byte3.cgate0.nand0.OUT VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1228 VSS gt_re1.I gt_re1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1229 VSS a_145380_680# a_145340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1230 a_1060_190# a_120_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1231 byte4.buf_RE0.O byte4.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1232 a_53440_1090# a_52500_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1233 a_60720_190# byte3.dff_5.CLK a_60160_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1234 VDD gt_re3.I gt_re3.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1235 VSS a_123420_680# byte2.dff_5.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1236 VDD byte4.cgate0.latch0.I0.O byte4.cgate0.nand0.A VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1237 a_47640_1092# byte3.tinv1.ENB Do22 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1238 a_42100_190# a_41160_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1239 byte3.cgate0.latch0.I0.O byte3.cgate0.latch0.I0.ENB a_78600_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1240 VDD a_104520_680# a_104480_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1241 a_119040_190# byte2.dff_4.CLK a_118480_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1242 a_164070_190# byte1.dff_5.CLK a_163960_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1243 VSS a_156720_680# a_156680_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1244 a_4560_1090# a_4330_140# a_4000_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1245 VDD a_24060_680# a_24020_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1246 a_169500_306# byte1.tinv6.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1247 VDD a_44940_190# a_45600_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1248 VDD a_68880_680# a_68840_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1249 byte1.dff_2.O byte1.dff_2.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1250 Do2 byte1.tinv5.EN a_165720_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1251 VDD byte3.tinv4.I a_58980_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1252 a_78600_306# byte3.cgate0.latch0.I0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1253 VDD a_127200_680# a_127160_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1254 a_163680_1090# a_163450_140# a_163120_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1255 byte3.buf_RE0.O byte3.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1256 a_130980_680# a_130770_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1257 VDD byte4.buf_RE1.I byte4.buf_RE1.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1258 VSS a_56380_140# a_56280_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1259 VDD a_67620_190# a_68280_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1260 byte1.dff_0.O byte1.dff_0.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1261 VSS a_67720_140# a_67620_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1262 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1263 a_121080_306# byte2.tinv4.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1264 a_148950_190# a_148330_140# a_148840_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1265 VSS a_49980_680# byte3.dff_2.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1266 byte2.cgate0.latch0.I0.O byte2.cgate0.latch0.I0.O a_96420_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1267 a_163120_140# a_163450_140# a_163350_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1268 a_156120_1090# a_155890_140# a_155560_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1269 a_146820_1092# byte1.tinv0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1270 VDD byte1.inv_and.I byte1.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1271 byte4.buf_RE1.O byte4.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1272 a_49980_680# a_49770_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1273 VSS byte2.buf_RE0.I byte2.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1274 byte1.dff_6.O byte1.dff_6.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1275 a_43860_1092# byte3.tinv0.ENB Do23 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1276 byte2.dff_4.O byte2.dff_4.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1277 VSS byte1.buf_RE1.I byte1.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1278 a_160460_190# a_159670_140# a_160290_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1279 a_159570_1090# Di3 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1280 a_148000_140# byte1.dff_1.CLK a_148230_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1281 a_93000_306# byte2.nand.B VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1282 a_169500_1092# byte1.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1283 VSS byte1.tinv2.I a_154380_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1284 a_42100_1090# a_41160_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1285 a_64270_140# byte3.dff_6.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1286 a_150600_306# byte1.tinv1.EN Do6 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1287 VSS a_127200_680# a_127160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1288 byte2.dff_7.O byte2.dff_7.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1289 a_37200_1092# byte4.cgate0.latch0.I0.O byte4.cgate0.latch0.I0.O VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1290 a_78600_1092# byte3.cgate0.latch0.I0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1291 VSS a_57540_680# byte3.dff_4.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1292 VSS byte3.cgate0.nand0.A a_78240_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1293 a_152900_1090# byte1.dff_2.CLK a_152730_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1294 VDD a_41260_140# a_41160_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1295 VDD byte1.tinv4.I a_161940_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1296 VDD a_57540_680# a_57500_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1297 VSS a_68880_680# byte3.dff_7.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1298 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1299 a_52830_190# Di20 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1300 a_104520_680# a_104310_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1301 a_105960_306# byte2.tinv0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1302 byte2.dff_6.O byte2.dff_6.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1303 byte3.buf_RE1.O byte3.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1304 VDD a_170580_190# a_171240_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1305 gt_re2.O gt_re2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1306 a_114930_1090# Di12 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1307 VSS byte4.buf_RE0.I byte4.buf_RE0.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1308 a_103360_140# byte2.dff_0.CLK a_103590_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1309 byte2.buf_RE1.O byte2.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1310 a_145340_1090# byte1.dff_0.CLK a_145170_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1311 a_27520_1090# a_26580_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1312 VDD byte4.buf_RE0.I byte4.buf_RE0.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1313 byte3.cgate0.inv1.O byte3.cgate0.nand0.OUT VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1314 VSS buf_ck1.I buf_ck1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1315 a_107980_1090# a_107040_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1316 VDD a_115860_680# byte2.dff_3.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1317 byte4.dff_5.O byte4.dff_5.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1318 VSS a_42420_680# a_42380_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1319 VSS byte1.buf_RE0.I byte1.buf_RE0.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1320 VSS a_125940_190# a_126600_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1321 a_130940_190# a_130150_140# a_130770_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1322 VDD a_26680_140# a_26580_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1323 a_55200_306# byte3.tinv3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1324 a_108090_190# byte2.dff_1.CLK a_107980_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1325 a_111250_140# byte2.dff_2.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1326 a_126040_140# byte2.dff_6.CLK a_126270_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1327 VSS byte2.tinv5.I a_124860_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1328 Do7 byte1.tinv0.ENB a_146820_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1329 VDD byte1.cgate0.nand0.B byte1.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1330 byte4.dff_0.O byte4.dff_0.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1331 VDD a_19020_190# a_19680_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1332 a_60490_140# byte3.dff_5.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1333 byte2.cgate0.nand0.A byte2.cgate0.latch0.I0.O VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1334 buf_sel1.O buf_sel1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1335 Do21 byte3.tinv2.EN a_51420_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1336 VDD a_1380_680# a_1340_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1337 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1338 VDD byte2.cgate0.nand0.OUT byte2.cgate0.inv1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1339 a_122590_140# byte2.dff_5.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1340 byte4.cgate0.nand0.OUT byte4.cgate0.nand0.A a_34860_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1341 Do18 byte3.tinv5.EN a_62760_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1342 VDD a_129820_140# a_129720_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1343 a_130940_1090# byte2.dff_7.CLK a_130770_190# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1344 byte3.dff_3.O byte3.dff_3.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1345 byte3.cgate0.nand0.A byte3.cgate0.latch0.I0.O VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1346 a_169500_1092# byte1.tinv6.ENB Do1 VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1347 VSS a_155560_140# a_155460_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1348 a_158160_1092# byte1.tinv3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1349 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1350 byte2.dff_4.O byte2.dff_4.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1351 VDD byte3.cgate0.nand0.B byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1352 VSS a_166900_140# a_166800_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1353 a_16500_680# a_16290_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1354 byte3.buf_RE1.O byte3.buf_RE1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1355 gt_re1.O gt_re1.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1356 VSS a_41160_190# a_41820_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1357 a_130380_1090# a_130150_140# a_129820_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1358 a_15670_140# byte4.dff_4.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1359 VDD WE3 byte4.nand.OUT VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1360 VDD a_46200_680# a_46160_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1361 VDD a_112080_680# byte2.dff_2.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1362 Do28 byte4.tinv3.EN a_14160_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1363 a_24060_680# a_23850_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1364 byte2.dff_2.O byte2.dff_2.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1365 a_107140_140# a_107470_140# a_107370_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1366 VSS a_26580_190# a_27240_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1367 VDD a_22900_140# a_22800_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1368 a_103590_1090# Di15 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1369 VSS byte2.inv_and.I byte2.inv_and.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1370 a_118480_140# a_118810_140# a_118710_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1371 a_23130_1090# Di25 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1372 byte2.buf_RE0.O byte2.buf_RE0.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1373 a_113520_1092# byte2.tinv2.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1374 a_115650_190# a_115030_140# a_115540_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1375 a_118810_140# byte2.dff_4.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1376 a_130380_190# byte2.dff_7.CLK a_129820_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1377 byte1.buf_RE1.O byte1.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1378 VSS a_7680_190# a_8340_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1379 VSS gt_re3.I gt_re3.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1380 a_104480_190# a_103690_140# a_104310_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1381 a_127200_680# a_126990_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1382 a_16180_1090# a_15240_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1383 a_67950_1090# Di16 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1384 VDD a_104520_680# byte2.dff_0.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1385 a_23230_140# byte4.dff_6.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1386 a_126270_1090# Di9 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1387 VSS a_156720_680# byte1.dff_3.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1388 VDD a_15340_140# a_15240_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1389 a_114700_140# byte2.dff_3.CLK a_114930_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1390 VDD byte1.cgate0.latch0.I0.I a_136020_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1391 a_4330_140# byte4.dff_1.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1392 a_67720_140# a_68050_140# a_67950_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1393 a_105960_306# byte2.tinv0.EN Do15 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1394 a_152010_190# Di5 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1395 VDD a_120_190# a_780_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1396 a_45370_140# byte3.dff_1.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1397 VDD a_127200_680# byte2.dff_6.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1398 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1399 byte3.dff_2.O byte3.dff_2.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1400 a_56710_140# byte3.dff_4.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1401 a_78600_1092# byte3.cgate0.latch0.I0.ENB byte3.cgate0.latch0.I0.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1402 a_65060_190# a_64270_140# a_64890_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1403 VSS a_126040_140# a_125940_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1404 a_11890_140# byte4.dff_3.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1405 VSS byte3.tinv4.I a_58980_306# VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1406 byte2.buf_RE0.O byte2.buf_RE0.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1407 byte2.cgate0.latch0.I0.O byte2.cgate0.latch0.I0.O a_95160_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1408 a_164280_680# a_164070_190# VSS VSS nfet_03v3 ad=425f pd=2.7u as=425f ps=2.7u w=850n l=300n
X1409 a_55200_306# byte3.tinv3.EN Do20 VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1410 a_60720_1090# a_60490_140# a_60160_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1411 VDD byte3.inv_and.I byte3.inv_and.O VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1412 a_103920_190# byte2.dff_0.CLK a_103360_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1413 a_19120_140# a_19450_140# a_19350_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1414 a_23740_190# a_22800_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1415 a_111870_190# a_111250_140# a_111760_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1416 a_154380_306# byte1.tinv2.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1417 Do11 byte2.tinv4.ENB a_121080_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1418 a_4840_1090# a_3900_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1419 VDD buf_ck1.I buf_ck1.O VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1420 a_4840_190# a_3900_190# VSS VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1421 a_12720_680# a_12510_190# VDD VDD pfet_03v3 ad=850f pd=4.4u as=850f ps=4.4u w=1.7u l=300n
X1422 VDD a_20280_680# byte4.dff_5.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1423 a_52600_140# byte3.dff_3.CLK a_52830_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1424 Do6 byte1.tinv1.EN a_150600_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1425 a_220_140# a_550_140# a_450_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=212.5f ps=1.35u w=850n l=300n
X1426 a_16460_190# a_15670_140# a_16290_190# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1427 a_78240_306# byte3.cgate0.nand0.B byte3.cgate0.latch0.I0.O VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1428 VDD a_65100_680# byte3.dff_6.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1429 Do3 byte1.tinv4.EN a_161940_306# VSS nfet_03v3 ad=255f pd=1.45u as=510f ps=2.9u w=850n l=300n
X1430 byte1.dff_2.O byte1.dff_2.O_bar VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1431 byte3.dff_6.O byte3.dff_6.O_bar VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1432 byte2.buf_RE1.O byte2.buf_RE1.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1433 a_104310_190# a_103690_140# a_104200_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=212.5f ps=1.95u w=1.7u l=300n
X1434 a_167850_190# byte1.dff_6.CLK a_167740_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1435 a_27010_140# byte4.dff_7.CLK VDD VDD pfet_03v3 ad=850f pd=4.4u as=467.5f ps=2.25u w=1.7u l=300n
X1436 VSS a_41260_140# a_41160_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1437 gt_re3.O gt_re3.I VSS VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1438 Do13 byte2.tinv2.ENB a_113520_1092# VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1439 VSS a_149160_680# a_149120_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=106.25f ps=1.1u w=850n l=300n
X1440 a_56610_1090# Di19 VDD VDD pfet_03v3 ad=425f pd=2.2u as=467.5f ps=2.25u w=1.7u l=300n
X1441 a_64500_190# byte3.dff_6.CLK a_63940_140# VSS nfet_03v3 ad=106.25f pd=1.1u as=233.75f ps=1.4u w=850n l=300n
X1442 a_45040_140# byte3.dff_1.CLK a_45270_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1443 VSS a_52600_140# a_52500_190# VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1444 a_66540_1092# byte3.tinv6.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1445 VSS byte3.buf_RE1.I byte3.buf_RE1.O VSS nfet_03v3 ad=510f pd=2.9u as=255f ps=1.45u w=850n l=300n
X1446 VSS gt_re2.I gt_re2.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1447 a_111150_190# Di13 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1448 VDD byte1.tinv0.I a_146820_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1449 VSS a_127200_680# byte2.dff_6.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
X1450 a_49660_1090# a_48720_190# VDD VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1451 VSS byte2.buf_RE1.I byte2.buf_RE1.O VSS nfet_03v3 ad=255f pd=1.45u as=255f ps=1.45u w=850n l=300n
X1452 a_171010_140# byte1.dff_7.CLK VSS VSS nfet_03v3 ad=425f pd=2.7u as=233.75f ps=1.4u w=850n l=300n
X1453 VDD a_57540_680# byte3.dff_4.O_bar VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1454 a_122490_190# Di10 VSS VSS nfet_03v3 ad=212.5f pd=1.35u as=233.75f ps=1.4u w=850n l=300n
X1455 VDD a_48820_140# a_48720_190# VDD pfet_03v3 ad=467.5f pd=2.25u as=850f ps=4.4u w=1.7u l=300n
X1456 a_119040_1090# a_118810_140# a_118480_140# VDD pfet_03v3 ad=212.5f pd=1.95u as=467.5f ps=2.25u w=1.7u l=300n
X1457 a_67720_140# byte3.dff_7.CLK a_67950_1090# VDD pfet_03v3 ad=467.5f pd=2.25u as=425f ps=2.2u w=1.7u l=300n
X1458 gt_re3.O gt_re3.I VDD VDD pfet_03v3 ad=510f pd=2.3u as=510f ps=2.3u w=1.7u l=300n
X1459 VDD byte1.tinv6.I a_169500_1092# VDD pfet_03v3 ad=1.02p pd=4.6u as=510f ps=2.3u w=1.7u l=300n
X1460 byte1.cgate0.nand0.OUT byte1.cgate0.nand0.A VDD VDD pfet_03v3 ad=510f pd=2.3u as=1.02p ps=4.6u w=1.7u l=300n
X1461 VSS a_20280_680# byte4.dff_5.O_bar VSS nfet_03v3 ad=233.75f pd=1.4u as=425f ps=2.7u w=850n l=300n
.ends

